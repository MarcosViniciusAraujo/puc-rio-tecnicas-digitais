CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 610 30 100 10
149 80 1278 651
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
317 176 430 273
42991634 0
0
6 Title:
5 Name:
0
0
0
44
13 Logic Switch~
5 509 433 0 1 11
0 27
0
0 0 21360 90
2 0V
14 0 28 8
3 V16
10 -10 31 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
331 0 0
2
5.90045e-315 0
0
13 Logic Switch~
5 734 438 0 10 11
0 35 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
14 0 28 8
3 V15
10 -10 31 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9604 0 0
2
5.90045e-315 0
0
13 Logic Switch~
5 679 437 0 1 11
0 34
0
0 0 21360 90
2 0V
14 0 28 8
3 V14
10 -10 31 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7518 0 0
2
5.90045e-315 0
0
13 Logic Switch~
5 544 433 0 10 11
0 28 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
14 0 28 8
3 V13
10 -10 31 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4832 0 0
2
5.90045e-315 0
0
13 Logic Switch~
5 630 435 0 1 11
0 33
0
0 0 21360 90
2 0V
14 0 28 8
3 V12
10 -10 31 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6798 0 0
2
5.90045e-315 0
0
13 Logic Switch~
5 582 433 0 1 11
0 32
0
0 0 21360 90
2 0V
14 0 28 8
3 V11
10 -10 31 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3336 0 0
2
5.90045e-315 0
0
13 Logic Switch~
5 11 98 0 1 11
0 36
0
0 0 21360 270
2 0V
-6 -21 8 -13
3 V10
-10 -31 11 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8370 0 0
2
5.90045e-315 0
0
13 Logic Switch~
5 16 354 0 1 11
0 37
0
0 0 21360 90
2 0V
11 0 25 8
2 V9
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3910 0 0
2
5.90045e-315 0
0
13 Logic Switch~
5 204 359 0 1 11
0 42
0
0 0 21360 90
2 0V
11 0 25 8
2 V8
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
316 0 0
2
5.90045e-315 0
0
13 Logic Switch~
5 150 359 0 1 11
0 41
0
0 0 21360 90
2 0V
11 0 25 8
2 V7
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
536 0 0
2
5.90045e-315 0
0
13 Logic Switch~
5 93 359 0 1 11
0 40
0
0 0 21360 90
2 0V
11 0 25 8
2 V6
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4460 0 0
2
5.90045e-315 0
0
13 Logic Switch~
5 49 354 0 10 11
0 39 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V5
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3260 0 0
2
5.90045e-315 0
0
13 Logic Switch~
5 53 111 0 10 11
0 43 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5156 0 0
2
5.90045e-315 0
0
13 Logic Switch~
5 100 111 0 1 11
0 44
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3133 0 0
2
5.90045e-315 0
0
13 Logic Switch~
5 135 114 0 1 11
0 45
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5523 0 0
2
5.90045e-315 0
0
13 Logic Switch~
5 171 113 0 1 11
0 46
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3746 0 0
2
5.90045e-315 0
0
7 Ground~
168 822 928 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5668 0 0
2
44816 0
0
7 Ground~
168 986 699 0 1 3
0 2
0
0 0 53360 180
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5368 0 0
2
44816 0
0
12 Hex Display~
7 904 1003 0 18 19
10 4 3 47 48 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 0 0 0 0
4 DISP
8293 0 0
2
44816 0
0
12 Hex Display~
7 966 1005 0 18 19
10 8 7 6 5 0 0 0 0 0
0 1 0 1 1 1 1 1 6
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
3232 0 0
2
44816 0
0
8 Hex Key~
166 758 985 0 11 12
0 12 11 10 9 0 0 0 0 0
6 54
0
0 0 4656 692
0
4 KPD1
19 -2 47 6
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
6644 0 0
2
44816 0
0
7 74LS283
152 1066 788 0 14 29
0 2 2 13 14 2 2 2 2 15
49 50 3 4 51
0
0 0 4848 0
6 74F283
-21 -60 21 -52
2 U8
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 14 3 5 11 15 2 6 7
10 13 1 4 9 12 14 3 5 11
15 2 6 7 10 13 1 4 9 0
65 0 0 512 0 0 0 0
1 U
4978 0 0
2
44816 0
0
7 74LS283
152 873 835 0 14 29
0 16 17 18 19 9 10 11 12 2
5 6 7 8 15
0
0 0 4848 0
6 74F283
-21 -60 21 -52
2 U7
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 14 3 5 11 15 2 6 7
10 13 1 4 9 12 14 3 5 11
15 2 6 7 10 13 1 4 9 0
65 0 0 0 0 0 0 0
1 U
9207 0 0
2
44816 0
0
5 4081~
219 404 614 0 3 22
0 20 26 13
0
0 0 624 270
4 4081
-7 -24 21 -16
3 U6B
16 -4 37 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 2 0
1 U
6998 0 0
2
44816 0
0
5 4081~
219 482 613 0 3 22
0 21 26 14
0
0 0 624 270
4 4081
-7 -24 21 -16
3 U6A
16 -4 37 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
3175 0 0
2
44816 0
0
5 4081~
219 547 612 0 3 22
0 22 26 16
0
0 0 624 270
4 4081
-7 -24 21 -16
3 U5D
16 -4 37 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 1 0
1 U
3378 0 0
2
44816 0
0
5 4081~
219 617 611 0 3 22
0 23 26 17
0
0 0 624 270
4 4081
-7 -24 21 -16
3 U5C
16 -4 37 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 1 0
1 U
922 0 0
2
44816 0
0
5 4081~
219 683 609 0 3 22
0 24 26 18
0
0 0 624 270
4 4081
-7 -24 21 -16
3 U5B
16 -4 37 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 1 0
1 U
6891 0 0
2
44816 0
0
5 4081~
219 749 609 0 3 22
0 25 26 19
0
0 0 624 270
4 4081
-7 -24 21 -16
3 U5A
16 -4 37 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
5407 0 0
2
44816 0
0
14 Logic Display~
6 389 42 0 1 2
10 20
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7349 0 0
2
5.90045e-315 0
0
14 Logic Display~
6 422 42 0 1 2
10 21
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3919 0 0
2
5.90045e-315 0
0
14 Logic Display~
6 449 43 0 1 2
10 22
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9747 0 0
2
5.90045e-315 0
0
14 Logic Display~
6 475 43 0 1 2
10 23
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5310 0 0
2
5.90045e-315 0
0
14 Logic Display~
6 500 44 0 1 2
10 24
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4318 0 0
2
5.90045e-315 0
0
14 Logic Display~
6 526 44 0 1 2
10 25
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3917 0 0
2
5.90045e-315 0
0
7 Ground~
168 851 135 0 1 3
0 2
0
0 0 53360 90
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7930 0 0
2
5.90045e-315 0
0
7 Ground~
168 1013 344 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6128 0 0
2
5.90045e-315 0
0
14 Logic Display~
6 1065 408 0 1 2
10 26
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L6
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7346 0 0
2
5.90045e-315 0
0
6 74LS85
106 904 265 0 14 29
0 2 2 20 21 2 2 27 28 31
30 29 26 52 53
0
0 0 5104 512
5 74F85
-18 -52 17 -44
2 U4
-7 -62 7 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 1 0 0 0
1 U
8577 0 0
2
5.90045e-315 0
0
6 74LS85
106 739 267 0 14 29
0 22 23 24 25 32 33 34 35 2
2 2 31 30 29
0
0 0 5104 0
5 74F85
-18 -52 17 -44
2 U3
-7 -62 7 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 0 1 0 0 0
1 U
3372 0 0
2
5.90045e-315 0
0
7 Ground~
168 211 481 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3741 0 0
2
5.90045e-315 0
0
4 4008
219 353 422 0 14 29
0 2 2 2 37 2 2 2 36 38
21 20 54 55 56
0
0 0 4848 0
4 4008
-14 -60 14 -52
2 U2
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
5813 0 0
2
5.90045e-315 0
0
7 Ground~
168 250 274 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3213 0 0
2
5.90045e-315 0
0
4 4008
219 269 205 0 14 29
0 43 44 45 46 39 40 41 42 2
25 24 23 22 38
0
0 0 4848 0
4 4008
-14 -60 14 -52
2 U1
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 0 1 0 0 0
1 U
3694 0 0
2
5.90045e-315 0
0
85
2 12 3 0 0 12432 0 19 22 0 0 5
907 1027
907 1056
1106 1056
1106 797
1098 797
13 1 4 0 0 8320 0 22 19 0 0 5
1098 806
1102 806
1102 1068
913 1068
913 1027
10 4 5 0 0 8320 0 23 20 0 0 5
905 826
940 826
940 1042
957 1042
957 1029
11 3 6 0 0 8320 0 23 20 0 0 5
905 835
945 835
945 1037
963 1037
963 1029
12 2 7 0 0 8320 0 23 20 0 0 5
905 844
993 844
993 1042
969 1042
969 1029
13 1 8 0 0 8320 0 23 20 0 0 5
905 853
988 853
988 1037
975 1037
975 1029
1 9 2 0 0 4096 0 17 23 0 0 3
822 922
822 880
841 880
0 8 2 0 0 0 0 0 22 9 0 3
1026 805
1026 815
1034 815
0 7 2 0 0 0 0 0 22 10 0 3
1026 796
1026 806
1034 806
0 6 2 0 0 0 0 0 22 11 0 4
986 787
1026 787
1026 797
1034 797
0 5 2 0 0 8192 0 0 22 12 0 3
986 751
986 788
1034 788
0 2 2 0 0 0 0 0 22 13 0 4
986 751
1026 751
1026 761
1034 761
1 1 2 0 0 0 0 18 22 0 0 3
986 707
986 752
1034 752
4 5 9 0 0 4224 0 21 23 0 0 3
749 961
749 835
841 835
3 6 10 0 0 4224 0 21 23 0 0 3
755 961
755 844
841 844
2 7 11 0 0 4224 0 21 23 0 0 3
761 961
761 853
841 853
1 8 12 0 0 4224 0 21 23 0 0 3
767 961
767 862
841 862
3 3 13 0 0 4224 0 22 24 0 0 3
1034 770
402 770
402 637
3 4 14 0 0 8320 0 25 22 0 0 3
480 636
480 779
1034 779
14 9 15 0 0 4224 0 23 22 0 0 4
905 880
1011 880
1011 833
1034 833
3 1 16 0 0 8320 0 26 23 0 0 3
545 635
545 799
841 799
3 2 17 0 0 8320 0 27 23 0 0 3
615 634
615 808
841 808
3 3 18 0 0 4224 0 28 23 0 0 3
681 632
681 817
841 817
3 4 19 0 0 4224 0 29 23 0 0 3
747 632
747 826
841 826
1 0 20 0 0 4096 0 24 0 0 39 4
411 592
411 427
389 427
389 422
1 0 21 0 0 4096 0 25 0 0 43 2
489 591
489 154
1 0 22 0 0 12416 0 26 0 0 61 4
554 590
554 448
468 448
468 185
0 1 23 0 0 4224 0 0 27 62 0 2
624 195
624 589
0 1 24 0 0 4224 0 0 28 63 0 2
690 205
690 587
0 1 25 0 0 4096 0 0 29 64 0 4
655 214
655 462
756 462
756 587
2 0 26 0 0 4096 0 28 0 0 35 2
672 587
672 481
2 0 26 0 0 4096 0 27 0 0 35 2
606 589
606 481
2 0 26 0 0 4096 0 26 0 0 35 2
536 590
536 481
2 0 26 0 0 4096 0 25 0 0 35 2
471 591
471 481
0 2 26 0 0 4224 0 0 24 36 0 3
739 481
393 481
393 592
0 2 26 0 0 0 0 0 29 37 0 4
868 412
868 481
738 481
738 587
12 1 26 0 0 0 0 39 38 0 0 4
872 283
868 283
868 412
1049 412
0 3 20 0 0 4224 0 0 39 39 0 4
389 122
991 122
991 256
936 256
11 1 20 0 0 0 0 42 30 0 0 3
385 422
389 422
389 60
1 7 27 0 0 8320 0 1 39 0 0 5
510 420
510 328
949 328
949 292
936 292
0 1 22 0 0 0 0 0 32 76 0 3
468 129
449 129
449 61
0 1 23 0 0 0 0 0 33 75 0 5
513 102
492 102
492 76
475 76
475 61
0 4 21 0 0 4224 0 0 39 44 0 4
413 154
949 154
949 265
936 265
10 1 21 0 0 0 0 42 31 0 0 5
385 431
413 431
413 115
422 115
422 60
1 0 2 0 0 4096 0 42 0 0 68 3
321 386
224 386
224 440
0 11 2 0 0 0 0 0 40 47 0 3
779 249
779 258
771 258
0 10 2 0 0 0 0 0 40 48 0 3
779 240
779 249
771 249
1 9 2 0 0 8192 0 36 40 0 0 4
844 136
779 136
779 240
771 240
0 1 2 0 0 0 0 0 39 52 0 4
1013 293
1014 293
1014 238
936 238
0 2 2 0 0 0 0 0 39 52 0 3
1007 292
1007 247
936 247
0 5 2 0 0 0 0 0 39 52 0 3
975 292
975 274
936 274
6 1 2 0 0 0 0 39 37 0 0 5
936 283
954 283
954 292
1013 292
1013 338
1 8 28 0 0 8320 0 4 39 0 0 5
545 420
545 323
944 323
944 301
936 301
14 11 29 0 0 4224 0 40 39 0 0 4
771 303
854 303
854 256
872 256
13 10 30 0 0 4224 0 40 39 0 0 4
771 294
859 294
859 247
872 247
12 9 31 0 0 4224 0 40 39 0 0 4
771 285
864 285
864 238
872 238
1 5 32 0 0 4224 0 6 40 0 0 3
583 420
583 276
707 276
1 6 33 0 0 4224 0 5 40 0 0 3
631 422
631 285
707 285
1 7 34 0 0 4224 0 3 40 0 0 3
680 424
680 294
707 294
1 8 35 0 0 4224 0 2 40 0 0 5
735 425
735 317
699 317
699 303
707 303
0 1 22 0 0 128 0 0 40 76 0 4
468 185
684 185
684 240
707 240
0 2 23 0 0 0 0 0 40 75 0 4
506 195
689 195
689 249
707 249
0 3 24 0 0 0 0 0 40 74 0 4
536 205
694 205
694 258
707 258
0 4 25 0 0 0 0 0 40 73 0 4
574 214
699 214
699 267
707 267
2 0 2 0 0 0 0 42 0 0 68 3
321 395
247 395
247 440
3 0 2 0 0 0 0 42 0 0 68 3
321 404
267 404
267 440
5 0 2 0 0 0 0 42 0 0 68 3
321 422
292 422
292 440
0 6 2 0 0 0 0 0 42 69 0 4
211 440
313 440
313 431
321 431
1 7 2 0 0 8320 0 41 42 0 0 3
211 475
211 440
321 440
1 8 36 0 0 20608 0 7 42 0 0 6
11 110
10 110
10 333
-1 333
-1 449
321 449
1 4 37 0 0 16512 0 8 42 0 0 5
17 341
17 338
2 338
2 413
321 413
14 9 38 0 0 8320 0 44 42 0 0 6
301 169
311 169
311 355
259 355
259 458
321 458
1 10 25 0 0 16512 0 35 44 0 0 5
526 62
526 95
574 95
574 214
301 214
1 11 24 0 0 128 0 34 44 0 0 6
500 62
519 62
519 179
536 179
536 205
301 205
0 12 23 0 0 128 0 0 44 0 0 5
513 95
513 178
506 178
506 196
301 196
13 0 22 0 0 0 0 44 0 0 0 3
301 187
468 187
468 125
9 1 2 0 0 0 0 44 43 0 0 5
237 241
233 241
233 260
250 260
250 268
1 5 39 0 0 8320 0 12 44 0 0 3
50 341
50 205
237 205
1 6 40 0 0 8320 0 11 44 0 0 3
94 346
94 214
237 214
1 7 41 0 0 4224 0 10 44 0 0 3
151 346
151 223
237 223
1 8 42 0 0 4224 0 9 44 0 0 3
205 346
205 232
237 232
1 1 43 0 0 8320 0 13 44 0 0 3
53 123
53 169
237 169
1 2 44 0 0 8320 0 14 44 0 0 3
100 123
100 178
237 178
1 3 45 0 0 8320 0 15 44 0 0 3
135 126
135 187
237 187
1 4 46 0 0 4224 0 16 44 0 0 3
171 125
171 196
237 196
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
