CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1278 651
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
5
7 Ground~
168 115 396 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
4299 0 0
2
44815.7 0
0
8 Hex Key~
166 58 107 0 11 12
0 20 3 22 21 0 0 0 0 0
0 48
0
0 0 4656 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
9672 0 0
2
44815.7 0
0
7 74LS139
118 212 259 0 14 29
0 21 22 2 27 28 29 23 24 25
26 30 31 32 33
0
0 0 4848 0
7 74LS139
-24 -51 25 -43
2 U3
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
113 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+[%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 13 14 15 7 6 5
4 9 10 11 12 3 2 1 13 14
15 7 6 5 4 9 10 11 12 0
65 0 0 512 0 0 0 0
1 U
7876 0 0
2
44815.7 0
0
7 74LS139
118 385 334 0 14 29
0 3 20 25 3 20 26 11 10 9
8 7 6 5 4
0
0 0 4848 0
7 74LS139
-24 -51 25 -43
2 U2
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
113 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+[%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 13 14 15 7 6 5
4 9 10 11 12 3 2 1 13 14
15 7 6 5 4 9 10 11 12 0
65 0 0 0 0 0 0 0
1 U
6369 0 0
2
44815.7 0
0
7 74LS139
118 385 201 0 14 29
0 3 20 23 3 20 24 12 13 14
15 16 17 18 19
0
0 0 4848 0
7 74LS139
-24 -51 25 -43
2 U1
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
113 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+[%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 13 14 15 7 6 5
4 9 10 11 12 3 2 1 13 14
15 7 6 5 4 9 10 11 12 0
65 0 0 0 0 0 0 0
1 U
9172 0 0
2
44815.7 0
0
31
0 2 3 0 0 4224 0 0 2 24 0 4
335 183
62 183
62 131
61 131
1 3 2 0 0 4224 0 1 3 0 0 3
115 390
115 259
174 259
0 14 4 0 0 4224 0 0 4 0 0 2
499 370
423 370
0 13 5 0 0 4224 0 0 4 0 0 2
499 361
423 361
0 12 6 0 0 4224 0 0 4 0 0 2
499 352
423 352
0 11 7 0 0 4224 0 0 4 0 0 2
499 343
423 343
0 10 8 0 0 4224 0 0 4 0 0 2
499 334
423 334
0 9 9 0 0 4224 0 0 4 0 0 2
499 325
423 325
0 8 10 0 0 4224 0 0 4 0 0 2
499 316
423 316
0 7 11 0 0 4224 0 0 4 0 0 2
499 307
423 307
7 0 12 0 0 4224 0 5 0 0 0 2
423 174
499 174
8 0 13 0 0 4224 0 5 0 0 0 2
423 183
499 183
9 0 14 0 0 4224 0 5 0 0 0 2
423 192
499 192
10 0 15 0 0 4224 0 5 0 0 0 2
423 201
499 201
11 0 16 0 0 4224 0 5 0 0 0 2
423 210
499 210
12 0 17 0 0 4224 0 5 0 0 0 2
423 219
499 219
13 0 18 0 0 4224 0 5 0 0 0 2
423 228
499 228
14 0 19 0 0 4224 0 5 0 0 0 2
423 237
499 237
0 4 3 0 0 0 0 0 4 21 0 4
329 315
314 315
314 352
353 352
0 5 20 0 0 8192 0 0 4 22 0 4
323 325
339 325
339 361
353 361
0 1 3 0 0 0 0 0 4 24 0 4
335 219
329 219
329 316
353 316
0 2 20 0 0 8192 0 0 4 23 0 4
322 226
323 226
323 325
353 325
0 5 20 0 0 0 0 0 5 25 0 3
322 192
322 228
353 228
4 1 3 0 0 128 0 5 5 0 0 4
353 219
335 219
335 183
353 183
1 2 20 0 0 12432 0 2 5 0 0 4
67 131
77 131
77 192
353 192
4 1 21 0 0 8320 0 2 3 0 0 3
49 131
49 241
180 241
3 2 22 0 0 8320 0 2 3 0 0 3
55 131
55 250
180 250
7 3 23 0 0 4224 0 3 5 0 0 4
250 232
339 232
339 201
347 201
8 6 24 0 0 4224 0 3 5 0 0 4
250 241
339 241
339 237
347 237
9 3 25 0 0 4224 0 3 4 0 0 4
250 250
334 250
334 334
347 334
10 6 26 0 0 8320 0 3 4 0 0 4
250 259
319 259
319 370
347 370
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
