CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1278 651
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
10
13 Logic Switch~
5 108 507 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V2
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.90046e-315 0
0
13 Logic Switch~
5 65 508 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V1
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.90046e-315 0
0
12 Hex Display~
7 653 159 0 18 19
10 6 5 4 3 0 0 0 0 0
0 1 1 1 1 1 1 1 8
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3124 0 0
2
5.90046e-315 0
0
7 Ground~
168 337 574 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3421 0 0
2
5.90046e-315 0
0
8 Hex Key~
166 249 97 0 11 12
0 21 17 13 9 0 0 0 0 0
8 56
0
0 0 4656 0
0
4 KPD4
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
8157 0 0
2
5.90046e-315 0
0
8 Hex Key~
166 183 95 0 11 12
0 22 18 14 10 0 0 0 0 0
2 50
0
0 0 4656 0
0
4 KPD3
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
5572 0 0
2
5.90046e-315 0
0
8 Hex Key~
166 125 96 0 11 12
0 23 19 15 11 0 0 0 0 0
6 54
0
0 0 4656 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
8901 0 0
2
5.90046e-315 0
0
8 Hex Key~
166 65 96 0 11 12
0 24 20 16 12 0 0 0 0 0
2 50
0
0 0 4656 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
7361 0 0
2
5.90046e-315 0
0
4 4539
219 406 394 0 14 29
0 13 14 15 16 2 9 10 11 12
2 7 8 3 4
0
0 0 4848 0
4 4539
-14 -60 14 -52
2 U2
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 4 5 6 1 13 12 11 10
15 2 14 9 7 3 4 5 6 1
13 12 11 10 15 2 14 9 7 0
65 0 0 0 1 0 0 0
1 U
4747 0 0
2
5.90046e-315 0
0
4 4539
219 405 215 0 14 29
0 21 22 23 24 2 17 18 19 20
2 7 8 5 6
0
0 0 4848 0
4 4539
-14 -60 14 -52
2 U1
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 4 5 6 1 13 12 11 10
15 2 14 9 7 3 4 5 6 1
13 12 11 10 15 2 14 9 7 0
65 0 0 0 1 0 0 0
1 U
972 0 0
2
5.90046e-315 0
0
28
13 4 3 0 0 8320 0 9 3 0 0 3
438 421
644 421
644 183
14 3 4 0 0 4224 0 9 3 0 0 3
438 376
650 376
650 183
13 2 5 0 0 4224 0 10 3 0 0 3
437 242
656 242
656 183
14 1 6 0 0 4224 0 10 3 0 0 3
437 197
662 197
662 183
10 0 2 0 0 4096 0 9 0 0 8 4
368 439
342 439
342 440
337 440
5 0 2 0 0 4096 0 9 0 0 8 2
368 394
337 394
10 0 2 0 0 0 0 10 0 0 8 2
367 260
337 260
5 1 2 0 0 8320 0 10 4 0 0 3
367 215
337 215
337 568
0 11 7 0 0 4096 0 0 10 10 0 4
66 448
354 448
354 269
373 269
1 11 7 0 0 8320 0 2 9 0 0 3
66 495
66 448
374 448
0 12 8 0 0 4096 0 0 10 12 0 4
109 457
359 457
359 278
373 278
1 12 8 0 0 8320 0 1 9 0 0 3
109 494
109 457
374 457
6 4 9 0 0 8320 0 9 5 0 0 3
374 403
240 403
240 121
7 4 10 0 0 8320 0 9 6 0 0 3
374 412
174 412
174 119
8 4 11 0 0 8320 0 9 7 0 0 3
374 421
116 421
116 120
9 4 12 0 0 4224 0 9 8 0 0 3
374 430
56 430
56 120
3 1 13 0 0 4224 0 5 9 0 0 3
246 121
246 358
374 358
3 2 14 0 0 4224 0 6 9 0 0 3
180 119
180 367
374 367
3 3 15 0 0 4224 0 7 9 0 0 3
122 120
122 376
374 376
3 4 16 0 0 8320 0 8 9 0 0 3
62 120
62 385
374 385
2 6 17 0 0 8320 0 5 10 0 0 3
252 121
252 224
373 224
2 7 18 0 0 8320 0 6 10 0 0 3
186 119
186 233
373 233
2 8 19 0 0 8320 0 7 10 0 0 3
128 120
128 242
373 242
2 9 20 0 0 8320 0 8 10 0 0 3
68 120
68 251
373 251
1 1 21 0 0 8320 0 5 10 0 0 3
258 121
258 179
373 179
1 2 22 0 0 8320 0 6 10 0 0 3
192 119
192 188
373 188
1 3 23 0 0 8320 0 7 10 0 0 3
134 120
134 197
373 197
1 4 24 0 0 8320 0 8 10 0 0 3
74 120
74 206
373 206
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
