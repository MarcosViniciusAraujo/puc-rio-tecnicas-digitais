CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 100 10
176 80 1278 651
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
19
13 Logic Switch~
5 142 116 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.9005e-315 0
0
9 Inverter~
13 348 484 0 2 22
0 3 4
0
0 0 608 180
6 74LS04
-21 -19 21 -11
3 U4C
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 2 0
1 U
391 0 0
2
5.9005e-315 0
0
9 Inverter~
13 341 513 0 2 22
0 5 6
0
0 0 608 180
6 74LS04
-21 -19 21 -11
3 U4B
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
3124 0 0
2
5.9005e-315 0
0
5 4073~
219 282 433 0 4 22
0 17 6 4 14
0
0 0 608 90
4 4073
-7 -24 21 -16
3 U7B
16 -5 37 3
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 5 0
1 U
3421 0 0
2
5.9005e-315 0
0
8 2-In OR~
219 250 146 0 3 22
0 17 24 8
0
0 0 608 0
6 74LS32
-21 -24 21 -16
3 U8B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
8157 0 0
2
5.9005e-315 0
0
8 2-In OR~
219 243 247 0 3 22
0 18 24 7
0
0 0 608 0
6 74LS32
-21 -24 21 -16
3 U8A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
5572 0 0
2
5.9005e-315 0
0
9 2-In NOR~
219 317 348 0 3 22
0 14 13 9
0
0 0 608 90
6 74LS02
-21 -24 21 -16
3 U2A
31 0 52 8
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
8901 0 0
2
5.9005e-315 0
0
5 4073~
219 366 433 0 4 22
0 18 3 19 13
0
0 0 608 90
4 4073
-7 -24 21 -16
3 U7A
16 -5 37 3
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 5 0
1 U
7361 0 0
2
5.9005e-315 0
0
2 +V
167 521 512 0 1 3
0 20
0
0 0 54240 270
2 5V
-7 -15 7 -7
2 V4
-7 -25 7 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4747 0 0
2
5.9005e-315 0
0
5 4082~
219 464 481 0 5 22
0 20 10 11 12 19
0
0 0 608 180
4 4082
-7 -24 21 -16
3 U5A
-13 -28 8 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 3 0
1 U
972 0 0
2
5.9005e-315 0
0
12 Hex Display~
7 713 69 0 16 19
10 3 21 16 15 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3472 0 0
2
5.9005e-315 0
0
12 Hex Display~
7 759 70 0 18 19
10 12 11 10 5 0 0 0 0 0
0 0 0 1 1 1 1 1 11
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
9998 0 0
2
5.9005e-315 0
0
7 Ground~
168 536 294 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3536 0 0
2
5.9005e-315 0
0
9 Inverter~
13 180 202 0 2 22
0 17 18
0
0 0 608 270
6 74LS04
-21 -19 21 -11
3 U4A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
4597 0 0
2
5.9005e-315 0
0
7 Pulser~
4 133 173 0 10 12
0 26 27 24 28 0 0 5 5 4
7
0
0 0 4640 0
0
2 V3
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3835 0 0
2
5.9005e-315 0
0
7 74LS193
137 577 222 0 14 29
0 22 23 9 2 2 2 2 17 29
30 15 16 21 3
0
0 0 4832 0
6 74F193
-21 -51 21 -43
2 U3
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 5 4 11 14 9 10 1 15 12
13 7 6 2 3 5 4 11 14 9
10 1 15 12 13 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
3670 0 0
2
5.9005e-315 0
0
7 Ground~
168 328 225 0 1 3
0 2
0
0 0 53344 270
0
4 GND1
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5616 0 0
2
5.9005e-315 0
0
2 +V
167 331 263 0 1 3
0 25
0
0 0 54240 90
2 5V
-7 -15 7 -7
2 V1
-7 -25 7 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9323 0 0
2
5.9005e-315 0
0
7 74LS193
137 437 225 0 14 29
0 8 7 9 2 2 25 25 25 22
23 5 10 11 12
0
0 0 4832 0
6 74F193
-21 -51 21 -43
2 U1
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 5 4 11 14 9 10 1 15 12
13 7 6 2 3 5 4 11 14 9
10 1 15 12 13 7 6 2 3 0
65 0 0 0 1 0 0 0
1 U
317 0 0
2
5.9005e-315 0
0
45
1 0 3 0 0 4096 0 2 0 0 23 3
369 484
409 484
409 459
3 2 4 0 0 8320 0 4 2 0 0 3
290 454
290 484
333 484
1 0 5 0 0 8320 0 3 0 0 9 3
362 513
488 513
488 234
3 0 4 0 0 0 0 4 0 0 2 2
290 454
290 459
2 2 6 0 0 4224 0 4 3 0 0 3
281 454
281 513
326 513
2 3 7 0 0 4224 0 19 6 0 0 4
405 207
284 207
284 247
276 247
3 1 8 0 0 4224 0 5 19 0 0 4
283 146
391 146
391 198
405 198
3 0 9 0 0 0 0 7 0 0 16 2
323 315
323 315
11 4 5 0 0 0 0 19 12 0 0 5
469 234
515 234
515 102
750 102
750 94
0 3 10 0 0 4096 0 0 12 28 0 3
515 325
756 325
756 94
0 2 11 0 0 4224 0 0 12 29 0 3
510 338
762 338
762 94
0 1 12 0 0 4224 0 0 12 30 0 3
505 349
768 349
768 94
4 0 2 0 0 4096 0 16 0 0 32 3
545 222
545 231
537 231
4 0 2 0 0 4096 0 19 0 0 42 3
405 225
373 225
373 234
0 3 9 0 0 4224 0 0 16 16 0 4
323 306
522 306
522 213
539 213
0 3 9 0 0 0 0 0 19 0 0 5
323 319
323 268
386 268
386 216
399 216
4 2 13 0 0 8320 0 8 7 0 0 4
365 409
365 379
332 379
332 367
4 1 14 0 0 8320 0 4 7 0 0 4
281 409
281 379
314 379
314 367
11 4 15 0 0 8320 0 16 11 0 0 3
609 231
704 231
704 93
12 3 16 0 0 8320 0 16 11 0 0 3
609 240
710 240
710 93
0 1 17 0 0 4224 0 0 4 40 0 4
212 116
212 483
272 483
272 454
0 1 18 0 0 4224 0 0 8 37 0 4
183 237
183 463
356 463
356 454
2 0 3 0 0 8320 0 8 0 0 27 4
365 454
365 459
637 459
637 258
5 3 19 0 0 8320 0 10 8 0 0 4
437 481
437 495
374 495
374 454
1 1 20 0 0 4224 0 10 9 0 0 4
482 494
502 494
502 511
509 511
13 2 21 0 0 8320 0 16 11 0 0 3
609 249
716 249
716 93
14 1 3 0 0 0 0 16 11 0 0 3
609 258
722 258
722 93
12 2 10 0 0 8336 0 19 10 0 0 4
469 243
515 243
515 485
482 485
13 3 11 0 0 0 0 19 10 0 0 4
469 252
510 252
510 476
482 476
14 4 12 0 0 0 0 19 10 0 0 4
469 261
505 261
505 467
482 467
7 6 2 0 0 0 0 16 16 0 0 2
545 249
545 240
6 0 2 0 0 0 0 16 0 0 33 3
545 240
545 231
537 231
5 1 2 0 0 8192 0 16 13 0 0 3
545 231
536 231
536 288
0 8 17 0 0 0 0 0 16 40 0 4
230 116
518 116
518 258
545 258
9 1 22 0 0 4224 0 19 16 0 0 4
475 216
526 216
526 195
545 195
10 2 23 0 0 4224 0 19 16 0 0 4
475 225
531 225
531 204
545 204
2 1 18 0 0 0 0 14 6 0 0 3
183 220
183 238
230 238
2 0 24 0 0 8320 0 6 0 0 41 3
230 256
205 256
205 164
0 1 17 0 0 0 0 0 14 40 0 2
183 116
183 184
1 1 17 0 0 0 0 1 5 0 0 4
154 116
230 116
230 137
237 137
3 2 24 0 0 0 0 15 5 0 0 4
157 164
230 164
230 155
237 155
1 5 2 0 0 8320 0 17 19 0 0 3
335 226
335 234
405 234
0 6 25 0 0 8192 0 0 19 44 0 3
391 252
391 243
405 243
0 7 25 0 0 0 0 0 19 45 0 3
391 261
391 252
405 252
1 8 25 0 0 4224 0 18 19 0 0 2
342 261
405 261
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
