CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
170 390 30 110 10
176 80 1278 651
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.440191 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
46
13 Logic Switch~
5 57 1011 0 1 11
0 44
0
0 0 21360 0
2 0V
-6 -16 8 -8
4 INIC
-13 -26 15 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
44902.7 0
0
13 Logic Switch~
5 148 1071 0 10 11
0 34 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
5 CLOCK
-16 -26 19 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
44902.7 1
0
13 Logic Switch~
5 531 849 0 1 11
0 47
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
44902.7 2
0
8 2-In OR~
219 719 1058 0 3 22
0 3 4 5
0
0 0 624 180
6 74LS32
-21 -24 21 -16
4 U18C
-2 -25 26 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
3421 0 0
2
44902.7 0
0
8 2-In OR~
219 1086 916 0 3 22
0 9 10 7
0
0 0 624 90
6 74LS32
-21 -24 21 -16
4 U18B
29 -3 57 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
8157 0 0
2
44902.7 0
0
8 2-In OR~
219 390 716 0 3 22
0 6 11 12
0
0 0 624 90
6 74LS32
-21 -24 21 -16
4 U18A
29 -3 57 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
5572 0 0
2
44902.7 0
0
9 Inverter~
13 1084 780 0 2 22
0 7 13
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U13E
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 2 0
1 U
8901 0 0
2
44902.7 0
0
7 Ground~
168 1499 516 0 1 3
0 2
0
0 0 53360 0
0
5 GND12
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7361 0 0
2
44902.7 0
0
7 Ground~
168 1670 471 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
4747 0 0
2
44902.7 0
0
2 +V
167 1699 442 0 1 3
0 16
0
0 0 54256 270
2 5V
-7 -15 7 -7
2 V1
-7 -25 7 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
972 0 0
2
44902.7 0
0
7 74LS191
135 1623 404 0 14 29
0 2 6 8 2 2 2 2 16 93
94 17 18 19 20
0
0 0 4848 512
6 74F191
-21 -51 21 -43
3 U17
-11 -52 10 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 14 11 5 9 10 1 15 13
12 7 6 2 3 4 14 11 5 9
10 1 15 13 12 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
3472 0 0
2
44902.7 0
0
7 74LS157
122 1426 433 0 14 29
0 9 20 24 19 23 18 22 17 21
2 25 26 27 28
0
0 0 4848 512
6 74F157
-21 -60 21 -52
3 U16
-17 -61 4 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
9998 0 0
2
44902.7 0
0
9 Inverter~
13 337 1076 0 2 22
0 29 30
0
0 0 624 180
6 74LS04
-21 -19 21 -11
4 U13D
-8 -20 20 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 2 0
1 U
3536 0 0
2
44902.7 0
0
9 2-In AND~
219 397 1076 0 3 22
0 32 31 29
0
0 0 624 180
6 74LS08
-21 -24 21 -16
4 U14A
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
4597 0 0
2
44902.7 0
0
7 Ground~
168 446 1097 0 1 3
0 2
0
0 0 53360 180
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3835 0 0
2
44902.7 0
0
4 4028
219 511 1131 0 14 29
0 2 32 31 33 15 14 10 11 9
6 95 96 97 98
0
0 0 4848 0
4 4028
-14 -60 14 -52
3 U12
-11 -61 10 -53
0
15 DVDD=16;DGND=8;
106 %D [%16bi %8bi %1i %2i %3i %4i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 11 12 13 10 3 14 2 15 1
6 7 4 9 5 11 12 13 10 3
14 2 15 1 6 7 4 9 5 0
65 0 0 512 0 0 0 0
1 U
3670 0 0
2
44902.7 0
0
7 Ground~
168 278 1202 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5616 0 0
2
44902.7 0
0
7 74LS191
135 361 1140 0 14 29
0 5 34 30 2 2 2 2 2 99
100 101 32 31 33
0
0 0 4848 0
6 74F191
-21 -51 21 -43
3 U11
-10 -52 11 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 14 11 5 9 10 1 15 13
12 7 6 2 3 4 14 11 5 9
10 1 15 13 12 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
9323 0 0
2
44902.7 0
0
5 4082~
219 1120 675 0 5 22
0 35 36 37 38 3
0
0 0 624 270
4 4082
-7 -24 21 -16
4 U15A
20 -4 48 4
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 4 0
1 U
317 0 0
2
5.90057e-315 0
0
9 Inverter~
13 276 1011 0 2 22
0 44 8
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U13C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 2 0
1 U
3108 0 0
2
44902.7 6
0
12 Hex Display~
7 641 872 0 16 19
10 42 41 40 39 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
4299 0 0
2
44902.7 7
0
7 Ground~
168 1313 607 0 1 3
0 2
0
0 0 53360 0
0
5 GND11
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9672 0 0
2
44902.7 8
0
2 +V
167 1453 593 0 1 3
0 43
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V6
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7876 0 0
2
44902.7 9
0
7 Ground~
168 1140 594 0 1 3
0 2
0
0 0 53360 0
0
5 GND10
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6369 0 0
2
44902.7 10
0
7 Ground~
168 1043 637 0 1 3
0 2
0
0 0 53360 0
0
4 GND9
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9172 0 0
2
44902.7 11
0
7 Ground~
168 456 711 0 1 3
0 2
0
0 0 53360 0
0
4 GND8
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7100 0 0
2
44902.7 13
0
7 Ground~
168 434 358 0 1 3
0 2
0
0 0 53360 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3820 0 0
2
44902.7 14
0
7 Ground~
168 796 713 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7678 0 0
2
44902.7 16
0
7 Ground~
168 790 512 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
961 0 0
2
44902.7 17
0
2 +V
167 463 903 0 1 3
0 48
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3178 0 0
2
44902.7 24
0
7 74LS174
130 1393 586 0 14 29
0 14 2 2 28 27 26 25 43 102
103 21 22 23 24
0
0 0 4848 692
7 74LS174
-24 -51 25 -43
3 U10
-11 -53 10 -45
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 9 14 13 11 6 4 3 1 15
12 10 7 5 2 9 14 13 11 6
4 3 1 15 12 10 7 5 2 0
65 0 0 512 1 0 0 0
1 U
3409 0 0
2
44902.7 25
0
7 74LS245
64 1189 543 0 18 37
0 104 105 106 107 35 36 37 38 108
109 110 111 28 27 26 25 2 13
0
0 0 4848 692
7 74LS245
-24 -60 25 -52
2 U9
-7 -62 7 -54
0
16 DVCC=20;DGND=10;
192 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i]
+ [%20bi %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP14
37

0 9 8 7 6 5 4 3 2 11
12 13 14 15 16 17 18 19 1 9
8 7 6 5 4 3 2 11 12 13
14 15 16 17 18 19 1 0
65 0 0 512 1 0 0 0
1 U
3951 0 0
2
44902.7 26
0
7 Ground~
168 994 633 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8885 0 0
2
44902.7 27
0
6 1K RAM
79 1031 552 0 20 41
0 2 2 49 50 51 52 53 54 55
56 112 113 114 115 35 36 37 38 2
13
0
0 0 4848 692
5 RAM1K
-17 -19 18 -11
2 U8
-7 -71 7 -63
0
16 DVCC=22;DGND=11;
214 %D [%22bi %11bi  %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i %19i %20i]
+ [%22bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o  %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o] %M
0
12 type:digital
5 DIP22
41

0 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 0
65 0 0 512 1 0 0 0
1 U
3780 0 0
2
44902.7 28
0
7 74LS157
122 835 646 0 14 29
0 7 60 68 59 67 58 66 57 65
2 52 51 50 49
0
0 0 4848 0
6 74F157
-21 -60 21 -52
2 U7
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
9265 0 0
2
44902.7 29
0
7 74LS157
122 837 437 0 14 29
0 7 64 72 63 71 62 70 61 69
2 56 55 54 53
0
0 0 4848 0
6 74F157
-21 -60 21 -52
2 U6
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
9442 0 0
2
44902.7 30
0
7 74LS191
135 547 761 0 14 29
0 2 45 8 2 77 78 79 80 116
117 57 58 59 60
0
0 0 4848 0
6 74F191
-21 -51 21 -43
2 U4
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 14 11 5 9 10 1 15 13
12 7 6 2 3 4 14 11 5 9
10 1 15 13 12 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
9424 0 0
2
44902.7 31
0
7 74LS191
135 553 645 0 14 29
0 2 12 8 2 81 82 83 84 45
118 61 62 63 64
0
0 0 4848 0
6 74F191
-21 -51 21 -43
2 U3
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 14 11 5 9 10 1 15 13
12 7 6 2 3 4 14 11 5 9
10 1 15 13 12 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
9968 0 0
2
44902.7 32
0
7 74LS191
135 549 432 0 14 29
0 2 46 8 2 85 86 87 88 119
120 65 66 67 68
0
0 0 4848 0
6 74F191
-21 -51 21 -43
2 U2
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 14 11 5 9 10 1 15 13
12 7 6 2 3 4 14 11 5 9
10 1 15 13 12 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
9281 0 0
2
44902.7 33
0
7 74LS191
135 546 278 0 14 29
0 2 6 8 2 89 90 91 92 46
121 69 70 71 72
0
0 0 4848 0
6 74F191
-21 -51 21 -43
2 U1
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 14 11 5 9 10 1 15 13
12 7 6 2 3 4 14 11 5 9
10 1 15 13 12 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
8464 0 0
2
44902.7 34
0
7 74LS191
135 539 920 0 14 29
0 47 6 8 48 73 74 75 76 122
4 39 40 41 42
0
0 0 4848 0
6 74F191
-21 -51 21 -43
2 U5
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 14 11 5 9 10 1 15 13
12 7 6 2 3 4 14 11 5 9
10 1 15 13 12 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
7168 0 0
2
44902.7 35
0
8 Hex Key~
166 99 822 0 11 12
0 76 75 74 73 0 0 0 0 0
4 52
0
0 0 4656 0
0
2 NP
-7 -34 7 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3171 0 0
2
44902.7 36
0
8 Hex Key~
166 101 679 0 11 12
0 80 79 78 77 0 0 0 0 0
0 48
0
0 0 4656 0
0
4 EDF2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
4139 0 0
2
44902.7 37
0
8 Hex Key~
166 101 560 0 11 12
0 84 83 82 81 0 0 0 0 0
10 65
0
0 0 4656 0
0
4 EDF1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
6435 0 0
2
44902.7 38
0
8 Hex Key~
166 102 323 0 11 12
0 88 87 86 85 0 0 0 0 0
0 48
0
0 0 4656 0
0
4 EDI2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
5283 0 0
2
44902.7 39
0
8 Hex Key~
166 100 193 0 11 12
0 92 91 90 89 0 0 0 0 0
1 49
0
0 0 4656 0
0
4 EDI1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
6874 0 0
2
44902.7 40
0
185
5 1 3 0 0 8320 0 19 4 0 0 3
1118 698
1118 1067
738 1067
0 2 4 0 0 20608 0 0 4 47 0 7
576 920
576 874
621 874
621 901
760 901
760 1049
738 1049
3 1 5 0 0 8336 0 4 18 0 0 5
692 1058
692 1049
310 1049
310 1113
323 1113
2 0 6 0 0 20608 0 11 0 0 8 7
1655 386
1665 386
1665 461
1656 461
1656 1126
586 1126
586 1131
1 0 7 0 0 4096 0 35 0 0 84 2
803 610
757 610
0 2 6 0 0 0 0 0 41 8 0 3
493 811
493 902
507 902
0 2 6 0 0 128 0 0 40 8 0 4
384 746
495 746
495 260
514 260
10 1 6 0 0 0 0 16 6 0 0 5
543 1131
587 1131
587 811
384 811
384 732
3 0 8 0 0 4096 0 11 0 0 12 2
1661 395
1723 395
0 1 9 0 0 4096 0 0 5 13 0 2
1080 1140
1080 932
2 7 10 0 0 8320 0 5 16 0 0 3
1098 932
1098 1158
543 1158
0 0 8 0 0 8320 0 0 0 0 58 4
1723 386
1723 1029
408 1029
408 1011
9 1 9 0 0 4224 0 16 12 0 0 4
543 1140
1486 1140
1486 397
1452 397
2 8 11 0 0 4224 0 6 16 0 0 5
402 732
402 1040
551 1040
551 1149
543 1149
3 2 12 0 0 8320 0 6 38 0 0 3
393 686
393 627
521 627
1 3 7 0 0 8320 0 7 5 0 0 4
1087 798
1088 798
1088 886
1089 886
20 0 13 0 0 8320 0 34 0 0 66 4
1069 571
1083 571
1083 718
1085 718
6 1 14 0 0 4224 0 16 31 0 0 4
543 1167
1353 1167
1353 605
1361 605
5 0 15 0 0 4224 0 16 0 0 0 4
543 1176
575 1176
575 1175
583 1175
10 1 2 0 0 4096 0 12 8 0 0 3
1458 478
1499 478
1499 510
4 0 2 0 0 0 0 11 0 0 25 2
1655 404
1670 404
5 0 2 0 0 0 0 11 0 0 25 2
1655 413
1670 413
6 0 2 0 0 0 0 11 0 0 25 2
1655 422
1670 422
7 0 2 0 0 0 0 11 0 0 25 2
1655 431
1670 431
1 1 2 0 0 8320 0 11 9 0 0 3
1661 377
1670 377
1670 465
8 1 16 0 0 4224 0 11 10 0 0 4
1655 440
1680 440
1680 441
1687 441
11 8 17 0 0 4224 0 11 12 0 0 4
1591 413
1491 413
1491 460
1452 460
12 6 18 0 0 4224 0 11 12 0 0 4
1591 422
1486 422
1486 442
1452 442
13 4 19 0 0 4224 0 11 12 0 0 4
1591 431
1481 431
1481 424
1452 424
14 2 20 0 0 4224 0 11 12 0 0 4
1591 440
1476 440
1476 406
1452 406
11 9 21 0 0 8320 0 31 12 0 0 4
1425 578
1463 578
1463 469
1452 469
12 7 22 0 0 8320 0 31 12 0 0 4
1425 569
1476 569
1476 451
1452 451
13 5 23 0 0 8320 0 31 12 0 0 4
1425 560
1471 560
1471 433
1452 433
14 3 24 0 0 8320 0 31 12 0 0 4
1425 551
1466 551
1466 415
1452 415
11 0 25 0 0 4224 0 12 0 0 97 2
1388 415
1284 415
12 1 26 0 0 4224 0 12 0 0 97 2
1388 433
1284 433
13 2 27 0 0 4224 0 12 0 0 97 2
1388 451
1284 451
14 3 28 0 0 4224 0 12 0 0 97 2
1388 469
1284 469
1 3 29 0 0 4224 0 13 14 0 0 2
358 1076
370 1076
3 2 30 0 0 8320 0 18 13 0 0 4
323 1131
315 1131
315 1076
322 1076
0 2 31 0 0 4224 0 0 14 45 0 3
436 1167
436 1067
415 1067
0 1 32 0 0 4096 0 0 14 44 0 3
425 1158
425 1085
415 1085
1 1 2 0 0 0 0 15 16 0 0 3
446 1105
446 1149
479 1149
12 2 32 0 0 4224 0 18 16 0 0 2
393 1158
479 1158
13 3 31 0 0 0 0 18 16 0 0 2
393 1167
479 1167
14 4 33 0 0 4224 0 18 16 0 0 2
393 1176
479 1176
10 0 4 0 0 144 0 41 0 0 0 2
571 920
581 920
1 2 34 0 0 4224 0 2 18 0 0 4
160 1071
290 1071
290 1122
329 1122
4 0 2 0 0 0 0 18 0 0 51 4
329 1140
289 1140
289 1160
292 1160
5 0 2 0 0 0 0 18 0 0 51 3
329 1149
300 1149
300 1159
0 6 2 0 0 0 0 0 18 52 0 5
292 1168
292 1159
300 1159
300 1158
329 1158
7 0 2 0 0 0 0 18 0 0 53 6
329 1167
292 1167
292 1168
283 1168
283 1178
278 1178
1 8 2 0 0 0 0 17 18 0 0 3
278 1196
278 1176
329 1176
1 0 35 0 0 12288 0 19 0 0 98 4
1131 653
1131 606
1126 606
1126 526
2 0 36 0 0 4224 0 19 0 0 99 4
1122 653
1122 522
1123 522
1123 517
3 0 37 0 0 4224 0 19 0 0 100 2
1113 653
1113 508
4 0 38 0 0 4224 0 19 0 0 101 2
1104 653
1104 499
2 3 8 0 0 0 0 20 41 0 0 4
297 1011
421 1011
421 911
501 911
11 4 39 0 0 4224 0 41 21 0 0 3
571 929
632 929
632 896
12 3 40 0 0 4224 0 41 21 0 0 3
571 938
638 938
638 896
13 2 41 0 0 4224 0 41 21 0 0 3
571 947
644 947
644 896
14 1 42 0 0 4224 0 41 21 0 0 3
571 956
650 956
650 896
2 0 2 0 0 0 0 31 0 0 64 3
1361 596
1333 596
1333 587
3 1 2 0 0 0 0 31 22 0 0 3
1361 587
1313 587
1313 601
8 1 43 0 0 4224 0 31 23 0 0 3
1431 605
1453 605
1453 602
2 18 13 0 0 0 0 7 32 0 0 6
1087 762
1085 762
1085 718
1225 718
1225 571
1221 571
17 1 2 0 0 0 0 32 24 0 0 3
1151 571
1140 571
1140 588
19 1 2 0 0 0 0 34 25 0 0 5
1069 580
1073 580
1073 623
1043 623
1043 631
0 3 8 0 0 0 0 0 40 70 0 3
424 424
424 269
508 269
0 3 8 0 0 128 0 0 39 71 0 3
424 636
424 423
511 423
0 3 8 0 0 0 0 0 38 72 0 3
421 753
421 636
515 636
0 3 8 0 0 0 0 0 37 58 0 3
421 912
421 752
509 752
1 1 44 0 0 4224 0 1 20 0 0 2
69 1011
261 1011
1 0 2 0 0 0 0 39 0 0 80 4
511 405
483 405
483 406
478 406
1 0 2 0 0 0 0 40 0 0 81 4
508 251
503 251
503 278
500 278
1 0 2 0 0 0 0 37 0 0 78 2
509 734
470 734
1 0 2 0 0 0 0 38 0 0 79 3
515 618
467 618
467 645
4 0 2 0 0 0 0 37 0 0 79 4
515 761
470 761
470 689
456 689
4 1 2 0 0 0 0 38 26 0 0 3
521 645
456 645
456 705
0 4 2 0 0 0 0 0 39 81 0 3
478 366
478 432
517 432
1 4 2 0 0 128 0 27 40 0 0 9
434 352
434 344
447 344
447 362
457 362
457 366
500 366
500 278
514 278
10 1 2 0 0 0 0 35 28 0 0 5
797 691
788 691
788 699
796 699
796 707
10 1 2 0 0 0 0 36 29 0 0 3
799 482
790 482
790 506
0 1 7 0 0 8320 0 0 36 16 0 4
1088 878
757 878
757 401
805 401
9 2 45 0 0 12416 0 38 37 0 0 6
591 636
595 636
595 714
501 714
501 743
515 743
9 2 46 0 0 8320 0 40 39 0 0 6
584 269
591 269
591 385
503 385
503 414
517 414
1 1 47 0 0 8320 0 41 3 0 0 4
501 893
501 858
543 858
543 849
1 4 48 0 0 8320 0 30 41 0 0 3
463 912
463 920
507 920
4 3 28 0 0 0 0 31 0 0 97 2
1361 578
1284 578
5 2 27 0 0 0 0 31 0 0 97 2
1361 569
1284 569
6 1 26 0 0 0 0 31 0 0 97 2
1361 560
1284 560
7 0 25 0 0 0 0 31 0 0 97 2
1361 551
1284 551
13 3 28 0 0 0 0 32 0 0 97 2
1221 526
1284 526
14 2 27 0 0 0 0 32 0 0 97 2
1221 517
1284 517
15 1 26 0 0 0 0 32 0 0 97 2
1221 508
1284 508
16 0 25 0 0 0 0 32 0 0 97 2
1221 499
1284 499
-150640 0 1 0 0 4128 0 0 0 0 0 2
1284 371
1284 704
15 5 35 0 0 4224 0 34 32 0 0 2
1063 526
1157 526
16 6 36 0 0 0 0 34 32 0 0 2
1063 517
1157 517
17 7 37 0 0 0 0 34 32 0 0 2
1063 508
1157 508
18 8 38 0 0 0 0 34 32 0 0 2
1063 499
1157 499
0 1 2 0 0 0 0 0 33 104 0 3
991 580
994 580
994 627
14 3 49 0 0 8320 0 35 34 0 0 4
867 682
978 682
978 562
999 562
2 1 2 0 0 0 0 34 34 0 0 4
999 571
983 571
983 580
999 580
13 4 50 0 0 8320 0 35 34 0 0 4
867 664
969 664
969 553
999 553
12 5 51 0 0 8320 0 35 34 0 0 4
867 646
955 646
955 544
999 544
11 6 52 0 0 8320 0 35 34 0 0 4
867 628
943 628
943 535
999 535
14 7 53 0 0 4224 0 36 34 0 0 4
869 473
934 473
934 526
999 526
13 8 54 0 0 4224 0 36 34 0 0 4
869 455
952 455
952 517
999 517
12 9 55 0 0 4224 0 36 34 0 0 4
869 437
965 437
965 508
999 508
11 10 56 0 0 4224 0 36 34 0 0 4
869 419
977 419
977 499
999 499
8 -154809 57 0 0 12288 0 35 0 0 144 4
803 673
782 673
782 732
711 732
6 -154810 58 0 0 8192 0 35 0 0 144 4
803 655
769 655
769 719
711 719
4 -154811 59 0 0 4096 0 35 0 0 144 2
803 637
711 637
2 -154812 60 0 0 4096 0 35 0 0 144 2
803 619
711 619
8 -154813 61 0 0 4096 0 36 0 0 144 2
805 464
711 464
6 -154814 62 0 0 4096 0 36 0 0 144 2
805 446
711 446
4 -154815 63 0 0 4096 0 36 0 0 144 2
805 428
711 428
2 -154816 64 0 0 4096 0 36 0 0 144 2
805 410
711 410
9 -154489 65 0 0 4096 0 35 0 0 144 4
803 682
748 682
748 714
711 714
7 -154490 66 0 0 4096 0 35 0 0 144 4
803 664
729 664
729 697
711 697
5 -154491 67 0 0 4096 0 35 0 0 144 2
803 646
711 646
3 -154492 68 0 0 4096 0 35 0 0 144 2
803 628
711 628
9 -154493 69 0 0 4096 0 36 0 0 144 2
805 473
711 473
7 -154494 70 0 0 4096 0 36 0 0 144 2
805 455
711 455
5 -154495 71 0 0 4096 0 36 0 0 144 2
805 437
711 437
3 -154496 72 0 0 4096 0 36 0 0 144 2
805 419
711 419
11 -154809 57 0 0 4224 0 37 0 0 144 2
579 770
711 770
12 -154810 58 0 0 4224 0 37 0 0 144 2
579 779
711 779
13 -154811 59 0 0 4224 0 37 0 0 144 2
579 788
711 788
14 -154812 60 0 0 4224 0 37 0 0 144 2
579 797
711 797
11 -154813 61 0 0 4224 0 38 0 0 144 2
585 654
711 654
12 -154814 62 0 0 4224 0 38 0 0 144 2
585 663
711 663
13 -154815 63 0 0 4224 0 38 0 0 144 2
585 672
711 672
14 -154816 64 0 0 4224 0 38 0 0 144 2
585 681
711 681
11 -154489 65 0 0 4224 0 39 0 0 144 2
581 441
711 441
12 -154490 66 0 0 4224 0 39 0 0 144 2
581 450
711 450
13 -154491 67 0 0 4224 0 39 0 0 144 2
581 459
711 459
14 -154492 68 0 0 4224 0 39 0 0 144 2
581 468
711 468
11 -154493 69 0 0 4224 0 40 0 0 144 2
578 287
711 287
12 -154494 70 0 0 4224 0 40 0 0 144 2
578 296
711 296
13 -154495 71 0 0 4224 0 40 0 0 144 2
578 305
711 305
14 -154496 72 0 0 4224 0 40 0 0 144 2
578 314
711 314
-865999395 0 1 0 0 4128 0 0 0 0 0 2
711 152
711 968
5 -58172 73 0 0 4096 0 41 0 0 185 2
507 929
335 929
6 -58173 74 0 0 4096 0 41 0 0 185 2
507 938
335 938
7 -58174 75 0 0 4096 0 41 0 0 185 2
507 947
335 947
8 -58175 76 0 0 4096 0 41 0 0 185 2
507 956
335 956
5 -13052985 77 0 0 4096 0 37 0 0 185 2
515 770
335 770
6 -13052986 78 0 0 4096 0 37 0 0 185 2
515 779
335 779
7 -13052987 79 0 0 4096 0 37 0 0 185 2
515 788
335 788
8 -13052988 80 0 0 4096 0 37 0 0 185 2
515 797
335 797
5 -13052989 81 0 0 4096 0 38 0 0 185 2
521 654
335 654
6 -13052990 82 0 0 4096 0 38 0 0 185 2
521 663
335 663
7 -13052991 83 0 0 4096 0 38 0 0 185 2
521 672
335 672
8 -13052992 84 0 0 4096 0 38 0 0 185 2
521 681
335 681
5 -13052793 85 0 0 4096 0 39 0 0 185 2
517 441
335 441
6 -13052794 86 0 0 4096 0 39 0 0 185 2
517 450
335 450
7 -13052795 87 0 0 4096 0 39 0 0 185 2
517 459
335 459
8 -13052796 88 0 0 4096 0 39 0 0 185 2
517 468
335 468
5 -13052797 89 0 0 4096 0 40 0 0 185 2
514 287
335 287
6 -13052798 90 0 0 4096 0 40 0 0 185 2
514 296
335 296
7 -13052799 91 0 0 4096 0 40 0 0 185 2
514 305
335 305
8 -13052800 92 0 0 4096 0 40 0 0 185 2
514 314
335 314
4 -13052985 77 0 0 8320 0 43 0 0 185 3
92 703
92 744
335 744
3 -13052986 78 0 0 8320 0 43 0 0 185 3
98 703
98 733
335 733
2 -13052987 79 0 0 8320 0 43 0 0 185 3
104 703
104 724
335 724
1 -13052988 80 0 0 8320 0 43 0 0 185 3
110 703
110 714
335 714
4 -13052989 81 0 0 8320 0 44 0 0 185 3
92 584
92 629
335 629
3 -13052990 82 0 0 8320 0 44 0 0 185 3
98 584
98 618
335 618
2 -13052991 83 0 0 8320 0 44 0 0 185 3
104 584
104 607
335 607
1 -13052992 84 0 0 8320 0 44 0 0 185 3
110 584
110 597
335 597
4 -13052793 85 0 0 8320 0 45 0 0 185 3
93 347
93 394
335 394
3 -13052794 86 0 0 8320 0 45 0 0 185 3
99 347
99 379
335 379
2 -13052795 87 0 0 8320 0 45 0 0 185 3
105 347
105 367
335 367
1 -13052796 88 0 0 8320 0 45 0 0 185 3
111 347
111 356
335 356
4 -13052797 89 0 0 8320 0 46 0 0 185 3
91 217
91 251
335 251
3 -13052798 90 0 0 8320 0 46 0 0 185 3
97 217
97 241
335 241
2 -13052799 91 0 0 8320 0 46 0 0 185 3
103 217
103 233
335 233
1 -13052800 92 0 0 8320 0 46 0 0 185 3
109 217
109 225
335 225
4 -58172 73 0 0 8320 0 42 0 0 185 3
90 846
90 902
335 902
3 -58173 74 0 0 8320 0 42 0 0 185 3
96 846
96 897
335 897
2 -58174 75 0 0 8320 0 42 0 0 185 3
102 846
102 892
335 892
1 -58175 76 0 0 8320 0 42 0 0 185 3
108 846
108 888
335 888
-902506802 0 1 0 0 4256 0 0 0 0 0 2
335 144
335 963
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
