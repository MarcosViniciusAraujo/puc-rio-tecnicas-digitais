CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
60 0 30 110 10
176 80 1278 651
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
21
13 Logic Switch~
5 77 327 0 10 11
0 29 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
44822.8 0
0
7 Pulser~
4 673 387 0 10 12
0 30 31 32 3 0 0 5 5 2
8
0
0 0 4656 0
0
2 V3
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
391 0 0
2
44822.8 0
0
2 +V
167 791 407 0 1 3
0 4
0
0 0 54256 90
2 5V
-8 -15 6 -7
2 V2
-7 -25 7 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3124 0 0
2
5.90047e-315 0
0
14 Logic Display~
6 997 769 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3421 0 0
2
44822.8 1
0
5 4071~
219 727 899 0 3 22
0 9 5 8
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U6C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 3 0
1 U
8157 0 0
2
44822.8 2
0
14 Logic Display~
6 987 564 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5572 0 0
2
44822.8 3
0
5 4069~
219 647 594 0 2 22
0 14 12
0
0 0 624 0
4 4069
-7 -24 21 -16
3 U7A
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 1 4 0
1 U
8901 0 0
2
44822.8 4
0
5 4001~
219 798 636 0 3 22
0 9 13 15
0
0 0 624 0
4 4001
-14 -24 14 -16
3 U5C
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 3 2 0
1 U
7361 0 0
2
44822.8 5
0
14 Logic Display~
6 987 350 0 1 2
10 16
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4747 0 0
2
44822.8 6
0
14 Logic Display~
6 975 133 0 1 2
10 20
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
972 0 0
2
44822.8 7
0
5 4071~
219 797 486 0 3 22
0 18 9 17
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U6B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 3 0
1 U
3472 0 0
2
44822.8 8
0
5 4071~
219 821 243 0 3 22
0 9 23 22
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U6A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 3 0
1 U
9998 0 0
2
44822.8 9
0
5 4001~
219 875 884 0 3 22
0 10 8 7
0
0 0 624 0
4 4001
-14 -24 14 -16
3 U5B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 2 0
1 U
3536 0 0
2
44822.8 10
0
5 4001~
219 872 793 0 3 22
0 6 7 10
0
0 0 624 0
4 4001
-14 -24 14 -16
3 U5A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 2 0
1 U
4597 0 0
2
44822.8 11
0
6 74LS74
17 902 612 0 12 25
0 33 34 12 15 35 36 37 38 11
39 40 41
0
0 0 4848 0
6 74LS74
-21 -60 21 -52
2 U4
-7 -61 7 -53
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 3 2 4 1 11 12 10 13 5
6 9 8 3 2 4 1 11 12 10
13 5 6 9 8 0
65 0 0 512 1 0 0 0
1 U
3835 0 0
2
44822.8 12
0
6 74LS73
102 893 387 0 12 25
0 19 17 3 4 42 43 44 45 16
46 47 48
0
0 0 4848 0
6 74LS73
-21 -51 21 -43
2 U3
-7 -52 7 -44
0
15 DVCC=4;DGND=11;
111 %D [%4bi %11bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%4bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 14 3 1 2 7 10 5 6 12
13 9 8 14 3 1 2 7 10 5
6 12 13 9 8 0
65 0 0 512 1 0 0 0
1 U
3670 0 0
2
44822.8 13
0
5 4013~
219 888 194 0 6 22
0 21 49 50 22 51 20
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U2A
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 1 0
1 U
5616 0 0
2
44822.8 14
0
7 Ground~
168 380 361 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9323 0 0
2
44822.8 15
0
4 4514
219 418 260 0 30 45
0 25 26 27 28 24 2 9 21 23
19 18 14 13 6 5 52 53 54 55
56 57 58 0 0 0 0 0 0 0
4
0
0 0 4848 0
4 4514
-14 -87 14 -79
2 U1
-7 -88 7 -80
0
16 DVDD=24;DGND=12;
155 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 22 21 3 2 1 23 11 9 10
8 7 6 5 4 18 17 20 19 14
13 16 15 22 21 3 2 1 23 11
9 10 8 7 6 5 4 18 17 20
19 14 13 16 15 0
65 0 0 512 1 0 0 0
1 U
317 0 0
2
44822.8 16
0
14 NO PushButton~
191 135 322 0 2 5
0 24 29
0
0 0 4720 0
0
2 S2
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3108 0 0
2
44822.8 17
0
8 Hex Key~
166 123 175 0 11 12
0 28 27 26 25 0 0 0 0 0
4 52
0
0 0 4656 512
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
4299 0 0
2
44822.8 18
0
33
4 3 3 0 0 4224 0 2 16 0 0 4
703 387
837 387
837 378
855 378
1 4 4 0 0 4224 0 3 16 0 0 4
802 405
842 405
842 387
855 387
15 2 5 0 0 8320 0 19 5 0 0 4
450 260
508 260
508 908
714 908
14 1 6 0 0 8320 0 19 14 0 0 4
450 269
535 269
535 784
859 784
0 1 7 0 0 8320 0 0 4 8 0 3
923 884
997 884
997 787
3 2 8 0 0 4224 0 5 13 0 0 4
760 899
854 899
854 893
862 893
0 1 9 0 0 8192 0 0 5 15 0 4
738 626
706 626
706 890
714 890
3 2 7 0 0 0 0 13 14 0 0 6
914 884
923 884
923 813
851 813
851 802
859 802
3 1 10 0 0 8320 0 14 13 0 0 6
911 793
918 793
918 864
854 864
854 875
862 875
9 1 11 0 0 4224 0 15 6 0 0 3
934 585
987 585
987 582
2 3 12 0 0 4224 0 7 15 0 0 2
668 594
864 594
13 2 13 0 0 8320 0 19 8 0 0 4
450 278
591 278
591 645
785 645
12 1 14 0 0 8320 0 19 7 0 0 4
450 287
570 287
570 594
632 594
3 4 15 0 0 8320 0 8 15 0 0 4
837 636
856 636
856 603
864 603
0 1 9 0 0 0 0 0 8 18 0 3
738 495
738 627
785 627
9 1 16 0 0 4224 0 16 9 0 0 3
925 369
987 369
987 368
0 1 16 0 0 0 0 0 9 0 0 2
987 369
987 368
0 2 9 0 0 0 0 0 11 24 0 3
738 332
738 495
784 495
3 2 17 0 0 8320 0 11 16 0 0 4
830 486
847 486
847 369
861 369
11 1 18 0 0 4224 0 19 11 0 0 4
450 296
764 296
764 477
784 477
10 1 19 0 0 4224 0 19 16 0 0 4
450 305
847 305
847 360
861 360
6 1 20 0 0 4224 0 17 10 0 0 3
912 158
975 158
975 151
8 1 21 0 0 12416 0 19 17 0 0 5
450 323
487 323
487 129
888 129
888 137
7 1 9 0 0 4224 0 19 12 0 0 4
450 332
738 332
738 234
808 234
3 4 22 0 0 8320 0 12 17 0 0 3
854 243
888 243
888 200
9 2 23 0 0 4224 0 19 12 0 0 4
450 314
800 314
800 252
808 252
6 1 2 0 0 4224 0 19 18 0 0 2
380 287
380 355
1 5 24 0 0 4224 0 20 19 0 0 4
152 330
362 330
362 269
386 269
1 4 25 0 0 4224 0 19 21 0 0 3
386 215
132 215
132 199
3 2 26 0 0 8320 0 21 19 0 0 3
126 199
126 224
386 224
2 3 27 0 0 8320 0 21 19 0 0 3
120 199
120 233
386 233
1 4 28 0 0 8320 0 21 19 0 0 3
114 199
114 242
386 242
1 2 29 0 0 4224 0 1 20 0 0 4
89 327
110 327
110 330
118 330
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
