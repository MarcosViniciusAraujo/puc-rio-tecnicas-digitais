CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 1 100 10
176 80 1278 651
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
11
13 Logic Switch~
5 236 110 0 1 11
0 5
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.90048e-315 0
0
13 Logic Switch~
5 436 121 0 1 11
0 15
0
0 0 21360 180
2 0V
-7 -16 7 -8
2 V2
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
5.90048e-315 0
0
2 +V
167 548 91 0 1 3
0 3
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3124 0 0
2
5.90048e-315 0
0
12 Hex Display~
7 721 103 0 16 19
10 10 9 8 7 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3421 0 0
2
5.90048e-315 0
0
12 Hex Display~
7 767 103 0 16 19
10 14 13 12 11 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
8157 0 0
2
5.90048e-315 0
0
7 Ground~
168 415 179 0 1 3
0 2
0
0 0 53360 90
0
4 GND1
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5572 0 0
2
5.90048e-315 0
0
7 Pulser~
4 348 70 0 10 12
0 24 25 6 26 0 0 5 5 4
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
8901 0 0
2
5.90048e-315 0
0
8 Hex Key~
166 142 133 0 11 12
0 19 18 17 16 0 0 0 0 0
11 66
0
0 0 4656 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
7361 0 0
2
5.90048e-315 0
0
8 Hex Key~
166 179 133 0 11 12
0 23 22 21 20 0 0 0 0 0
13 68
0
0 0 4656 512
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
4747 0 0
2
5.90048e-315 0
0
7 74LS164
127 614 178 0 12 25
0 3 4 6 5 7 8 9 10 11
12 13 14
0
0 0 4848 0
6 74F164
-21 -51 21 -43
2 U2
-7 -52 7 -44
0
15 DVCC=14;DGND=7;
96 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 1 2 8 9 13 12 11 10 6
5 4 3 1 2 8 9 13 12 11
10 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
972 0 0
2
5.90048e-315 0
0
7 74LS165
97 305 198 0 14 29
0 16 17 18 19 20 21 22 23 15
5 2 6 27 4
0
0 0 4848 0
7 74LS165
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 6 5 4 3 14 13 12 11 10
1 15 2 7 9 6 5 4 3 14
13 12 11 10 1 15 2 7 9 0
65 0 0 512 1 0 0 0
1 U
3472 0 0
2
5.90048e-315 0
0
24
1 1 3 0 0 4224 0 3 10 0 0 3
548 100
548 151
582 151
14 2 4 0 0 4224 0 11 10 0 0 4
337 234
568 234
568 160
582 160
0 4 5 0 0 12416 0 0 10 13 0 4
356 141
361 141
361 196
576 196
0 3 6 0 0 4224 0 0 10 16 0 4
382 164
546 164
546 178
582 178
5 4 7 0 0 4224 0 10 4 0 0 3
646 151
712 151
712 127
6 3 8 0 0 4224 0 10 4 0 0 3
646 160
718 160
718 127
7 2 9 0 0 4224 0 10 4 0 0 3
646 169
724 169
724 127
8 1 10 0 0 4224 0 10 4 0 0 3
646 178
730 178
730 127
9 4 11 0 0 4224 0 10 5 0 0 3
646 187
758 187
758 127
10 3 12 0 0 4224 0 10 5 0 0 3
646 196
764 196
764 127
11 2 13 0 0 4224 0 10 5 0 0 3
646 205
770 205
770 127
12 1 14 0 0 4224 0 10 5 0 0 3
646 214
776 214
776 127
1 10 5 0 0 0 0 1 11 0 0 5
236 122
236 125
356 125
356 171
343 171
1 9 15 0 0 4224 0 2 11 0 0 4
422 121
351 121
351 162
337 162
11 1 2 0 0 4224 0 11 6 0 0 2
343 180
408 180
3 12 6 0 0 0 0 7 11 0 0 4
372 61
382 61
382 189
337 189
4 1 16 0 0 8320 0 8 11 0 0 3
133 157
133 171
273 171
3 2 17 0 0 8320 0 8 11 0 0 3
139 157
139 180
273 180
2 3 18 0 0 8320 0 8 11 0 0 3
145 157
145 189
273 189
1 4 19 0 0 8320 0 8 11 0 0 3
151 157
151 198
273 198
4 5 20 0 0 8320 0 9 11 0 0 3
188 157
188 207
273 207
3 6 21 0 0 8320 0 9 11 0 0 3
182 157
182 216
273 216
2 7 22 0 0 8320 0 9 11 0 0 3
176 157
176 225
273 225
1 8 23 0 0 8320 0 9 11 0 0 3
170 157
170 234
273 234
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
