CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 2030 30 100 10
176 80 1278 651
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
33
5 4082~
219 455 456 0 5 22
0 13 35 34 3 2
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U10B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 10 0
1 U
5130 0 0
2
44807.9 0
0
5 4049~
219 202 829 0 2 22
0 3 4
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U11B
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 11 0
1 U
391 0 0
2
44807.9 0
0
8 Hex Key~
166 76 43 0 11 12
0 3 11 12 13 0 0 0 0 0
8 56
0
0 0 4656 512
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
3124 0 0
2
44807.9 0
0
5 4071~
219 574 2485 0 3 22
0 7 6 5
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U6B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 6 0
1 U
3421 0 0
2
5.90045e-315 0
0
5 4049~
219 233 2648 0 2 22
0 3 8
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U11A
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 11 0
1 U
8157 0 0
2
5.90045e-315 0
0
5 4049~
219 238 2610 0 2 22
0 11 9
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U5F
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 5 0
1 U
5572 0 0
2
5.90045e-315 0
0
5 4049~
219 238 2573 0 2 22
0 12 10
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U5E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 5 0
1 U
8901 0 0
2
5.90045e-315 0
0
5 4082~
219 392 2605 0 5 22
0 13 10 9 8 6
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U10A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 10 0
1 U
7361 0 0
2
5.90045e-315 0
0
5 4069~
219 211 2361 0 2 22
0 12 14
0
0 0 624 0
4 4069
-7 -24 21 -16
3 U8C
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 3 8 0
1 U
4747 0 0
2
5.90045e-315 0
0
5 4069~
219 211 2323 0 2 22
0 13 15
0
0 0 624 0
4 4069
-7 -24 21 -16
3 U8B
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 2 8 0
1 U
972 0 0
2
5.90045e-315 0
0
5 4082~
219 377 2365 0 5 22
0 15 14 11 3 7
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U9B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 9 0
1 U
3472 0 0
2
5.90045e-315 0
0
8 3-In OR~
219 789 1709 0 4 22
0 19 18 17 16
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U3B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 3 0
1 U
9998 0 0
2
5.90045e-315 0
0
5 4049~
219 272 2001 0 2 22
0 3 20
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U5D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 5 0
1 U
3536 0 0
2
5.90045e-315 0
0
5 4049~
219 272 1830 0 2 22
0 13 21
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U5C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 5 0
1 U
4597 0 0
2
5.90045e-315 0
0
5 4082~
219 517 1920 0 5 22
0 21 12 11 20 17
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U9A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 9 0
1 U
3835 0 0
2
5.90045e-315 0
0
5 4069~
219 279 1709 0 2 22
0 11 22
0
0 0 624 0
4 4069
-7 -24 21 -16
3 U8A
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 1 8 0
1 U
3670 0 0
2
5.90045e-315 0
0
5 4069~
219 274 1639 0 2 22
0 12 23
0
0 0 624 0
4 4069
-7 -24 21 -16
3 U2F
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 6 2 0
1 U
5616 0 0
2
5.90045e-315 0
0
5 4073~
219 509 1709 0 4 22
0 23 22 3 18
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U7A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 7 0
1 U
9323 0 0
2
5.90045e-315 0
0
5 4069~
219 313 1466 0 2 22
0 11 24
0
0 0 624 0
4 4069
-7 -24 21 -16
3 U2E
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 5 2 0
1 U
317 0 0
2
5.90045e-315 0
0
5 4069~
219 316 1400 0 2 22
0 13 25
0
0 0 624 0
4 4069
-7 -24 21 -16
3 U2D
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 4 2 0
1 U
3108 0 0
2
5.90045e-315 0
0
5 4073~
219 497 1465 0 4 22
0 25 24 3 19
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U4C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 4 0
1 U
4299 0 0
2
5.90045e-315 0
0
5 4071~
219 663 850 0 3 22
0 28 27 26
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U6A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 6 0
1 U
9672 0 0
2
44807.9 0
0
5 4049~
219 186 995 0 2 22
0 11 29
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U5B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 5 0
1 U
7876 0 0
2
44807.9 1
0
5 4073~
219 461 950 0 4 22
0 30 12 29 27
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 4 0
1 U
6369 0 0
2
44807.9 2
0
5 4049~
219 260 735 0 2 22
0 13 30
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U5A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 5 0
1 U
9172 0 0
2
44807.9 3
0
5 4073~
219 454 777 0 4 22
0 30 11 4 28
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 4 0
1 U
7100 0 0
2
44807.9 4
0
12 Hex Display~
7 1029 74 0 18 19
10 31 26 16 5 0 0 0 0 0
0 1 1 1 1 1 1 1 8
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3820 0 0
2
44807.9 5
0
8 3-In OR~
219 653 310 0 4 22
0 33 32 2 31
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U3A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 3 0
1 U
7678 0 0
2
44807.9 6
0
5 4069~
219 253 474 0 2 22
0 12 35
0
0 0 624 0
4 4069
-7 -24 21 -16
3 U2C
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 3 2 0
1 U
961 0 0
2
44807.9 7
0
5 4069~
219 258 338 0 2 22
0 11 34
0
0 0 624 0
4 4069
-7 -24 21 -16
3 U2B
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 2 2 0
1 U
3178 0 0
2
44807.9 9
0
5 4073~
219 442 310 0 4 22
0 36 12 34 32
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 1 0
1 U
3409 0 0
2
44807.9 10
0
5 4069~
219 252 155 0 2 22
0 13 36
0
0 0 624 0
4 4069
-7 -24 21 -16
3 U2A
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 1 2 0
1 U
3951 0 0
2
44807.9 11
0
5 4073~
219 439 214 0 4 22
0 36 11 3 33
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 1 0
1 U
8885 0 0
2
44807.9 12
0
65
5 3 2 0 0 4224 0 1 28 0 0 4
476 456
632 456
632 319
640 319
0 4 3 0 0 4096 0 0 1 50 0 4
67 490
423 490
423 470
431 470
2 3 4 0 0 4224 0 2 26 0 0 3
223 829
430 829
430 786
3 4 5 0 0 8320 0 4 27 0 0 3
607 2485
1020 2485
1020 98
5 2 6 0 0 4224 0 8 4 0 0 4
413 2605
553 2605
553 2494
561 2494
5 1 7 0 0 4224 0 11 4 0 0 4
398 2365
553 2365
553 2476
561 2476
2 4 8 0 0 4224 0 5 8 0 0 3
254 2648
368 2648
368 2619
2 3 9 0 0 4224 0 6 8 0 0 2
259 2610
368 2610
2 2 10 0 0 4224 0 7 8 0 0 4
259 2573
356 2573
356 2601
368 2601
0 1 3 0 0 0 0 0 5 19 0 3
68 2431
68 2648
218 2648
0 1 11 0 0 4096 0 0 6 18 0 3
74 2391
74 2610
223 2610
0 1 12 0 0 4096 0 0 7 16 0 3
80 2361
80 2573
223 2573
0 1 13 0 0 8192 0 0 8 17 0 4
86 2322
86 2549
368 2549
368 2592
2 2 14 0 0 4224 0 9 11 0 0 2
232 2361
353 2361
2 1 15 0 0 4224 0 10 11 0 0 3
232 2323
353 2323
353 2352
0 1 12 0 0 4096 0 0 9 28 0 3
80 1888
80 2361
196 2361
0 1 13 0 0 4096 0 0 10 29 0 3
86 1828
86 2323
196 2323
0 3 11 0 0 4096 0 0 11 27 0 5
74 1955
74 2392
330 2392
330 2370
353 2370
0 4 3 0 0 4096 0 0 11 26 0 4
68 1999
68 2431
353 2431
353 2379
3 4 16 0 0 4224 0 27 12 0 0 3
1026 98
1026 1709
822 1709
5 3 17 0 0 4224 0 15 12 0 0 4
538 1920
762 1920
762 1718
776 1718
4 2 18 0 0 4224 0 18 12 0 0 2
530 1709
777 1709
4 1 19 0 0 4224 0 21 12 0 0 4
518 1465
767 1465
767 1700
776 1700
2 4 20 0 0 4224 0 13 15 0 0 4
293 2001
491 2001
491 1934
493 1934
2 1 21 0 0 4224 0 14 15 0 0 3
293 1830
493 1830
493 1907
0 1 3 0 0 0 0 0 13 32 0 4
67 1762
68 1762
68 2001
257 2001
0 3 11 0 0 0 0 0 15 33 0 6
73 1708
74 1708
74 1955
479 1955
479 1925
493 1925
0 2 12 0 0 0 0 0 15 39 0 6
79 1639
80 1639
80 1888
481 1888
481 1916
493 1916
0 1 13 0 0 0 0 0 14 36 0 3
86 1398
86 1830
257 1830
2 2 22 0 0 4224 0 16 18 0 0 2
300 1709
485 1709
2 1 23 0 0 4224 0 17 18 0 0 3
295 1639
485 1639
485 1700
0 3 3 0 0 0 0 0 18 37 0 4
67 1494
67 1766
485 1766
485 1718
0 1 11 0 0 0 0 0 16 38 0 3
73 1462
73 1709
264 1709
2 2 24 0 0 8320 0 19 21 0 0 3
334 1466
334 1465
473 1465
2 1 25 0 0 4224 0 20 21 0 0 3
337 1400
473 1400
473 1456
0 1 13 0 0 8320 0 0 20 47 0 4
85 735
86 735
86 1400
301 1400
0 3 3 0 0 4224 0 0 21 50 0 4
67 827
67 1496
473 1496
473 1474
0 1 11 0 0 4096 0 0 19 44 0 4
73 995
73 1465
298 1465
298 1466
0 1 12 0 0 4224 0 0 17 48 0 3
79 948
79 1639
259 1639
3 2 26 0 0 8320 0 22 27 0 0 3
696 850
1032 850
1032 98
4 2 27 0 0 4224 0 24 22 0 0 4
482 950
642 950
642 859
650 859
4 1 28 0 0 4224 0 26 22 0 0 4
475 777
642 777
642 841
650 841
2 3 29 0 0 4224 0 23 24 0 0 4
207 995
341 995
341 959
437 959
0 1 11 0 0 0 0 0 23 49 0 3
73 798
73 995
171 995
0 1 30 0 0 4224 0 0 24 46 0 3
307 735
307 941
437 941
2 1 30 0 0 0 0 25 26 0 0 4
281 735
422 735
422 768
430 768
0 1 13 0 0 0 0 0 25 57 0 3
85 441
85 735
245 735
0 2 12 0 0 0 0 0 24 60 0 3
79 310
79 950
437 950
0 2 11 0 0 4224 0 0 26 63 0 5
73 213
73 798
370 798
370 777
430 777
0 1 3 0 0 0 0 0 2 62 0 3
67 223
67 829
187 829
4 1 31 0 0 4224 0 28 27 0 0 3
686 310
1038 310
1038 98
4 2 32 0 0 4224 0 31 28 0 0 2
463 310
641 310
4 1 33 0 0 4224 0 33 28 0 0 4
460 214
632 214
632 301
640 301
0 3 34 0 0 4096 0 0 1 58 0 5
322 338
322 462
424 462
424 461
431 461
2 2 35 0 0 12416 0 29 1 0 0 4
274 474
315 474
315 452
431 452
0 1 12 0 0 0 0 0 29 60 0 3
143 310
143 474
238 474
0 1 13 0 0 0 0 0 1 65 0 3
85 155
85 443
431 443
2 3 34 0 0 4224 0 30 31 0 0 3
279 338
418 338
418 319
0 1 11 0 0 0 0 0 30 63 0 3
95 214
95 338
243 338
3 2 12 0 0 0 0 3 31 0 0 3
79 67
79 310
418 310
0 1 36 0 0 4224 0 0 31 64 0 3
310 155
310 301
418 301
1 3 3 0 0 0 0 3 33 0 0 3
67 67
67 223
415 223
2 2 11 0 0 0 0 3 33 0 0 3
73 67
73 214
415 214
2 1 36 0 0 0 0 32 33 0 0 4
273 155
407 155
407 205
415 205
4 1 13 0 0 0 0 3 32 0 0 3
85 67
85 155
237 155
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
