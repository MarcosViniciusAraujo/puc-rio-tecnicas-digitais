CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 30 30 70 10
176 80 1278 651
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
26
13 Logic Switch~
5 483 84 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
44857.9 0
0
13 Logic Switch~
5 451 84 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
391 0 0
2
44857.9 0
0
13 Logic Switch~
5 105 87 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 X0
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3124 0 0
2
44857.9 0
0
13 Logic Switch~
5 67 89 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 X1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3421 0 0
2
44857.9 0
0
9 Inverter~
13 704 117 0 2 22
0 4 3
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U4C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 6 0
1 U
8157 0 0
2
44857.9 0
0
14 Logic Display~
6 921 423 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5572 0 0
2
44857.9 0
0
5 4073~
219 783 460 0 4 22
0 11 10 9 8
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U8A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 10 0
1 U
8901 0 0
2
44857.9 0
0
5 4073~
219 239 785 0 4 22
0 15 14 13 12
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U3C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 5 0
1 U
7361 0 0
2
44857.9 0
0
5 4073~
219 235 693 0 4 22
0 13 16 14 18
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 5 0
1 U
4747 0 0
2
44857.9 0
0
5 4081~
219 237 633 0 3 22
0 13 10 19
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U6C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 8 0
1 U
972 0 0
2
44857.9 0
0
5 4081~
219 236 583 0 3 22
0 13 17 20
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U6B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 8 0
1 U
3472 0 0
2
44857.9 0
0
8 3-In OR~
219 394 628 0 4 22
0 20 19 18 21
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U7A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 9 0
1 U
9998 0 0
2
44857.9 0
0
5 4081~
219 229 351 0 3 22
0 9 14 22
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U6A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 8 0
1 U
3536 0 0
2
44857.9 0
0
5 4081~
219 222 407 0 3 22
0 15 9 23
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 4 0
1 U
4597 0 0
2
44857.9 0
0
5 4081~
219 231 466 0 3 22
0 13 24 25
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 4 0
1 U
3835 0 0
2
44857.9 0
0
5 4081~
219 228 516 0 3 22
0 15 14 26
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 4 0
1 U
3670 0 0
2
44857.9 0
0
8 4-In OR~
219 395 429 0 5 22
0 22 23 25 26 27
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U5A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 7 0
1 U
5616 0 0
2
44857.9 0
0
2 +V
167 466 278 0 1 3
0 28
0
0 0 54256 90
2 5V
-7 -15 7 -7
2 V1
-7 -25 7 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
9323 0 0
2
44857.9 0
0
9 Inverter~
13 77 139 0 2 22
0 14 17
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U4B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 6 0
1 U
317 0 0
2
44857.9 0
0
9 Inverter~
13 130 139 0 2 22
0 15 16
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U4A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 6 0
1 U
3108 0 0
2
44857.9 0
0
5 4073~
219 243 171 0 4 22
0 17 16 29 31
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 5 0
1 U
4299 0 0
2
44857.9 0
0
5 4081~
219 242 282 0 3 22
0 29 9 30
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 4 0
1 U
9672 0 0
2
44857.9 0
0
8 2-In OR~
219 389 238 0 3 22
0 31 30 32
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U1A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
7876 0 0
2
44857.9 0
0
5 4027~
219 538 679 0 7 32
0 5 21 7 12 3 9 24
0
0 0 4720 0
4 4027
7 -60 35 -52
2 Y2
25 -61 39 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 1 2 0
1 U
6369 0 0
2
44857.9 0
0
5 4027~
219 537 471 0 7 32
0 2 27 7 9 3 29 10
0
0 0 4720 0
4 4027
7 -60 35 -52
2 Y1
25 -61 39 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 2 1 0
1 U
9172 0 0
2
44857.9 0
0
5 4027~
219 534 294 0 7 32
0 33 32 7 28 3 11 13
0
0 0 4720 0
4 4027
7 -60 35 -52
2 Y0
21 -75 35 -67
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
7100 0 0
2
44857.9 0
0
51
0 5 3 0 0 4096 0 0 25 2 0 3
709 537
537 537
537 477
0 5 3 0 0 12416 0 0 24 3 0 6
707 359
707 308
709 308
709 693
538 693
538 685
2 5 3 0 0 16 0 5 26 0 0 4
707 135
707 359
534 359
534 300
1 1 4 0 0 8320 0 5 1 0 0 6
707 99
707 95
494 95
494 111
483 111
483 96
0 3 7 0 0 4224 0 0 24 6 0 3
451 444
451 652
514 652
0 3 7 0 0 0 0 0 25 7 0 3
451 289
451 444
513 444
3 1 7 0 0 0 0 26 2 0 0 4
510 267
510 289
451 289
451 96
4 1 8 0 0 4224 0 7 6 0 0 3
804 460
921 460
921 441
0 3 9 0 0 4096 0 0 7 47 0 2
591 469
759 469
0 2 10 0 0 4096 0 0 7 18 0 2
572 460
759 460
6 1 11 0 0 4224 0 26 7 0 0 4
564 276
751 276
751 451
759 451
4 4 12 0 0 4224 0 8 24 0 0 4
260 785
506 785
506 661
514 661
0 3 13 0 0 4096 0 0 8 35 0 3
49 457
49 794
215 794
0 2 14 0 0 8192 0 0 8 16 0 3
64 702
64 785
215 785
0 1 15 0 0 4096 0 0 8 36 0 3
104 507
104 776
215 776
0 3 14 0 0 8192 0 0 9 37 0 4
66 524
64 524
64 702
211 702
0 2 16 0 0 4224 0 0 9 43 0 3
133 171
133 693
211 693
7 2 10 0 0 12416 0 25 10 0 0 6
561 435
572 435
572 549
205 549
205 642
213 642
0 2 17 0 0 4224 0 0 11 42 0 3
80 160
80 592
212 592
0 1 13 0 0 0 0 0 9 21 0 4
143 624
142 624
142 684
211 684
0 1 13 0 0 0 0 0 10 22 0 3
143 572
143 624
213 624
0 1 13 0 0 0 0 0 11 35 0 3
143 457
143 574
212 574
4 3 18 0 0 4224 0 9 12 0 0 4
256 693
373 693
373 637
381 637
3 2 19 0 0 8320 0 10 12 0 0 3
258 633
258 628
382 628
3 1 20 0 0 4224 0 11 12 0 0 4
257 583
353 583
353 619
381 619
4 2 21 0 0 4224 0 12 24 0 0 4
427 628
506 628
506 643
514 643
0 2 9 0 0 0 0 0 14 28 0 3
188 340
188 416
198 416
0 1 9 0 0 0 0 0 13 47 0 3
188 318
188 342
205 342
0 2 14 0 0 0 0 0 13 37 0 2
66 360
205 360
0 1 15 0 0 0 0 0 14 36 0 4
104 399
119 399
119 398
198 398
1 3 22 0 0 4224 0 17 13 0 0 4
378 416
263 416
263 351
250 351
2 3 23 0 0 4224 0 17 14 0 0 4
378 425
259 425
259 407
243 407
0 4 9 0 0 0 0 0 25 47 0 3
591 499
513 499
513 453
7 2 24 0 0 12416 0 24 15 0 0 6
562 643
571 643
571 889
33 889
33 475
207 475
1 7 13 0 0 12416 0 15 26 0 0 6
207 457
34 457
34 50
572 50
572 258
558 258
0 1 15 0 0 8320 0 0 16 45 0 4
105 107
104 107
104 507
204 507
0 2 14 0 0 8320 0 0 16 46 0 4
67 108
66 108
66 525
204 525
3 3 25 0 0 4224 0 15 17 0 0 4
252 466
365 466
365 434
378 434
3 4 26 0 0 4224 0 16 17 0 0 4
249 516
370 516
370 443
378 443
5 2 27 0 0 4224 0 17 25 0 0 4
428 429
505 429
505 435
513 435
1 4 28 0 0 4224 0 18 26 0 0 2
477 276
510 276
2 1 17 0 0 0 0 19 21 0 0 3
80 157
80 162
219 162
2 2 16 0 0 0 0 20 21 0 0 3
133 157
133 171
219 171
3 0 29 0 0 8192 0 21 0 0 48 3
219 180
210 180
210 274
1 1 15 0 0 0 0 3 20 0 0 4
105 99
105 107
133 107
133 121
1 1 14 0 0 0 0 4 19 0 0 4
67 101
67 108
80 108
80 121
6 2 9 0 0 12416 0 24 22 0 0 6
568 661
591 661
591 318
175 318
175 291
218 291
6 1 29 0 0 12416 0 25 22 0 0 6
567 453
583 453
583 305
210 305
210 273
218 273
3 2 30 0 0 4224 0 22 23 0 0 4
263 282
368 282
368 247
376 247
4 1 31 0 0 4224 0 21 23 0 0 4
264 171
368 171
368 229
376 229
3 2 32 0 0 4224 0 23 26 0 0 4
422 238
508 238
508 258
510 258
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
