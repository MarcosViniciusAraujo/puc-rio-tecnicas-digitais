CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 630 4 100 10
176 80 1278 651
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
3 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
14
9 2-In AND~
219 267 937 0 3 22
0 4 3 6
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U2A
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
5130 0 0
2
5.90048e-315 0
0
7 Ground~
168 269 989 0 1 3
0 2
0
0 0 53360 270
0
4 GND2
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
391 0 0
2
5.90048e-315 0
0
7 Ground~
168 253 737 0 1 3
0 2
0
0 0 53360 270
0
4 GND1
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3124 0 0
2
5.90048e-315 0
0
6 74LS90
107 353 1021 0 10 21
0 2 2 6 6 7 5 18 19 4
5
0
0 0 4848 0
6 74LS90
-21 -51 21 -43
2 U3
-7 -52 7 -44
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 512 1 0 0 0
1 U
3421 0 0
2
5.90048e-315 0
0
7 Pulser~
4 173 873 0 10 12
0 20 21 8 22 0 0 5 5 5
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
8157 0 0
2
5.90048e-315 5.3568e-315
0
12 Hex Display~
7 640 785 0 18 19
10 3 9 10 7 0 0 0 0 0
0 1 0 1 1 0 1 1 5
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP4
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
5572 0 0
2
5.90048e-315 5.32571e-315
0
12 Hex Display~
7 587 783 0 16 19
10 5 4 23 24 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 1 0 0 0
4 DISP
8901 0 0
2
5.90048e-315 5.26354e-315
0
6 74LS90
107 358 779 0 10 21
0 2 2 6 6 8 3 7 10 9
3
0
0 0 4848 0
6 74LS90
-21 -51 21 -43
2 U1
-7 -52 7 -44
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 0 1 0 0 0
1 U
7361 0 0
2
5.90048e-315 0
0
5 4073~
219 264 489 0 4 22
0 12 16 15 11
0
0 0 624 180
4 4073
-7 -24 21 -16
3 U4B
-13 -25 8 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 2 0
1 U
4747 0 0
2
5.90048e-315 0
0
12 Hex Display~
7 584 335 0 16 19
10 12 25 26 27 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP3
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 1 0 0 0
4 DISP
972 0 0
2
5.90048e-315 0
0
6 74LS93
109 355 539 0 8 17
0 11 11 14 28 12 12 12 12
0
0 0 4848 0
6 74LS93
-21 -35 21 -27
2 U6
-7 -36 7 -28
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 512 1 0 0 0
1 U
3472 0 0
2
5.90048e-315 0
0
12 Hex Display~
7 637 337 0 18 19
10 16 13 15 14 0 0 0 0 0
0 1 0 1 1 0 1 1 5
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
9998 0 0
2
5.90048e-315 0
0
6 74LS93
109 355 413 0 8 17
0 11 11 17 16 14 15 13 16
0
0 0 4848 0
6 74LS93
-21 -35 21 -27
2 U5
-7 -36 7 -28
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 0 1 0 0 0
1 U
3536 0 0
2
5.90048e-315 0
0
7 Pulser~
4 170 425 0 10 12
0 29 30 17 31 0 0 5 5 5
7
0
0 0 4656 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
4597 0 0
2
5.90048e-315 0
0
39
0 2 3 0 0 8192 0 0 1 19 0 3
394 879
394 928
285 928
0 1 4 0 0 8192 0 0 1 3 0 3
411 1030
411 946
285 946
9 2 4 0 0 8320 0 4 7 0 0 3
385 1030
590 1030
590 807
6 0 5 0 0 12288 0 4 0 0 15 5
315 1048
311 1048
311 1068
414 1068
414 1048
0 2 2 0 0 8192 0 0 4 6 0 3
307 994
307 1003
321 1003
1 1 2 0 0 4096 0 2 4 0 0 4
276 990
307 990
307 994
321 994
2 0 2 0 0 0 0 8 0 0 8 4
326 761
315 761
315 752
312 752
1 1 2 0 0 4224 0 3 8 0 0 4
260 738
312 738
312 752
326 752
0 3 6 0 0 8192 0 0 4 10 0 3
307 1021
307 1012
321 1012
3 4 6 0 0 8192 0 1 4 0 0 4
240 937
237 937
237 1021
321 1021
5 0 7 0 0 16384 0 4 0 0 17 5
315 1039
307 1039
307 1090
436 1090
436 851
0 6 3 0 0 0 0 0 8 19 0 6
394 814
390 814
390 821
319 821
319 806
320 806
3 5 8 0 0 4224 0 5 8 0 0 4
197 864
312 864
312 797
320 797
4 0 6 0 0 0 0 8 0 0 20 3
326 779
326 770
317 770
10 1 5 0 0 8320 0 4 7 0 0 3
385 1048
596 1048
596 807
9 2 9 0 0 12416 0 8 6 0 0 5
390 788
408 788
408 870
643 870
643 809
7 4 7 0 0 12432 0 8 6 0 0 5
390 752
398 752
398 851
631 851
631 809
8 3 10 0 0 12416 0 8 6 0 0 5
390 770
403 770
403 861
637 861
637 809
10 1 3 0 0 20608 0 8 6 0 0 7
390 806
394 806
394 879
399 879
399 880
649 880
649 809
0 3 6 0 0 4224 0 0 8 10 0 3
238 937
238 770
326 770
0 2 11 0 0 8192 0 0 11 31 0 3
309 530
309 539
323 539
0 1 11 0 0 0 0 0 13 37 0 3
312 413
312 404
323 404
7 0 12 0 0 0 0 11 0 0 26 2
387 548
387 548
6 0 12 0 0 0 0 11 0 0 26 2
387 539
387 539
5 0 12 0 0 0 0 11 0 0 26 2
387 530
387 530
0 1 12 0 0 4224 0 0 10 32 0 3
391 557
593 557
593 359
7 2 13 0 0 4224 0 13 12 0 0 3
387 422
640 422
640 361
0 3 14 0 0 4096 0 0 11 33 0 5
433 404
433 572
309 572
309 548
317 548
0 3 15 0 0 8192 0 0 9 34 0 3
411 413
411 480
282 480
0 2 16 0 0 4096 0 0 9 38 0 3
315 454
315 489
282 489
4 1 11 0 0 12416 0 9 11 0 0 4
237 489
235 489
235 530
323 530
8 1 12 0 0 0 0 11 9 0 0 4
387 557
391 557
391 498
282 498
5 4 14 0 0 4224 0 13 12 0 0 3
387 404
628 404
628 361
6 3 15 0 0 4224 0 13 12 0 0 3
387 413
634 413
634 361
0 1 16 0 0 8320 0 0 12 38 0 4
396 431
396 432
646 432
646 361
0 3 17 0 0 0 0 0 13 39 0 2
317 422
317 422
0 2 11 0 0 0 0 0 13 31 0 3
235 489
235 413
323 413
8 4 16 0 0 0 0 13 13 0 0 6
387 431
396 431
396 454
314 454
314 431
317 431
3 3 17 0 0 4224 0 14 13 0 0 4
194 416
309 416
309 422
317 422
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
