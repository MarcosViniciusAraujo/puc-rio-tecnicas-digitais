CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1278 651
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
38
13 Logic Switch~
5 55 1624 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V10
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9281 0 0
2
44808.5 0
0
13 Logic Switch~
5 56 1572 0 1 11
0 7
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8464 0 0
2
44808.5 0
0
13 Logic Switch~
5 84 1223 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7168 0 0
2
44808.5 0
0
13 Logic Switch~
5 84 1165 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3171 0 0
2
44808.5 0
0
13 Logic Switch~
5 125 895 0 10 11
0 18 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4139 0 0
2
44808.4 0
0
13 Logic Switch~
5 125 843 0 1 11
0 17
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6435 0 0
2
44808.4 0
0
13 Logic Switch~
5 123 575 0 1 11
0 24
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
5283 0 0
2
44808.4 0
0
13 Logic Switch~
5 120 506 0 10 11
0 25 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
6874 0 0
2
44808.4 0
0
13 Logic Switch~
5 122 181 0 1 11
0 32
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
5305 0 0
2
44808.4 0
0
13 Logic Switch~
5 121 124 0 1 11
0 33
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
34 0 0
2
44808.4 0
0
14 Logic Display~
6 624 1617 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
969 0 0
2
44808.5 0
0
5 4030~
219 381 1644 0 3 22
0 4 5 3
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U6B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 6 0
1 U
8402 0 0
2
44808.5 0
0
5 4030~
219 163 1594 0 3 22
0 7 6 4
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U6A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 6 0
1 U
3751 0 0
2
44808.5 0
0
14 Logic Display~
6 599 1201 0 1 2
10 14
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4292 0 0
2
44808.5 0
0
5 4081~
219 391 1423 0 3 22
0 11 10 8
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U5D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 5 0
1 U
6118 0 0
2
44808.5 0
0
5 4081~
219 390 1336 0 3 22
0 13 12 9
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U5C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 5 0
1 U
34 0 0
2
44808.5 0
0
5 4030~
219 383 1229 0 3 22
0 12 13 14
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U4D
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 4 0
1 U
6357 0 0
2
44808.5 0
0
5 4030~
219 190 1193 0 3 22
0 10 11 12
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U4C
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 4 0
1 U
319 0 0
2
44808.5 0
0
5 4071~
219 524 1374 0 3 22
0 9 8 5
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U3D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 3 0
1 U
3976 0 0
2
44808.5 0
0
5 4071~
219 526 1000 0 3 22
0 16 15 13
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U3C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 3 0
1 U
7634 0 0
2
44808.4 0
0
5 4081~
219 399 1043 0 3 22
0 18 17 15
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 5 0
1 U
523 0 0
2
44808.4 0
0
5 4081~
219 398 969 0 3 22
0 19 20 16
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 5 0
1 U
6748 0 0
2
44808.4 0
0
14 Logic Display~
6 659 846 0 1 2
10 21
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6901 0 0
2
44808.4 0
0
5 4030~
219 384 871 0 3 22
0 20 19 21
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U4B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 4 0
1 U
842 0 0
2
44808.4 0
0
5 4030~
219 216 862 0 3 22
0 17 18 20
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U4A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 4 0
1 U
3277 0 0
2
44808.4 0
0
5 4071~
219 555 700 0 3 22
0 23 22 19
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 3 0
1 U
4212 0 0
2
44808.4 0
0
5 4081~
219 431 742 0 3 22
0 25 24 22
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 2 0
1 U
4720 0 0
2
44808.4 0
0
5 4081~
219 430 664 0 3 22
0 27 26 23
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 2 0
1 U
5551 0 0
2
44808.4 0
0
14 Logic Display~
6 648 529 0 1 2
10 28
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6986 0 0
2
44808.4 0
0
5 4030~
219 403 550 0 3 22
0 27 26 28
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U1D
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 1 0
1 U
8745 0 0
2
44808.4 0
0
5 4030~
219 231 541 0 3 22
0 25 24 27
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U1C
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 1 0
1 U
9592 0 0
2
44808.4 0
0
14 Logic Display~
6 642 170 0 1 2
10 29
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8748 0 0
2
44808.4 0
0
7 Ground~
168 67 265 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7168 0 0
2
44808.4 0
0
5 4071~
219 517 305 0 3 22
0 31 30 26
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 3 0
1 U
631 0 0
2
44808.4 0
0
5 4081~
219 410 349 0 3 22
0 33 32 30
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 2 0
1 U
9466 0 0
2
44808.4 0
0
5 4081~
219 408 278 0 3 22
0 34 2 31
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
3266 0 0
2
44808.4 0
0
5 4030~
219 397 191 0 3 22
0 34 2 29
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U1B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 1 0
1 U
7693 0 0
2
44808.4 0
0
5 4030~
219 241 143 0 3 22
0 33 32 34
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U1A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
3723 0 0
2
44808.4 0
0
49
3 1 3 0 0 4224 0 12 11 0 0 3
414 1644
624 1644
624 1635
1 3 4 0 0 4224 0 12 13 0 0 4
365 1635
204 1635
204 1594
196 1594
3 2 5 0 0 12432 0 19 12 0 0 6
557 1374
561 1374
561 1560
264 1560
264 1653
365 1653
1 2 6 0 0 4224 0 1 13 0 0 4
67 1624
137 1624
137 1603
147 1603
1 1 7 0 0 4224 0 2 13 0 0 4
68 1572
137 1572
137 1585
147 1585
3 2 8 0 0 4224 0 15 19 0 0 4
412 1423
503 1423
503 1383
511 1383
3 1 9 0 0 4224 0 16 19 0 0 4
411 1336
503 1336
503 1365
511 1365
2 0 10 0 0 8320 0 15 0 0 16 3
367 1432
104 1432
104 1165
1 0 11 0 0 4224 0 15 0 0 15 3
367 1414
140 1414
140 1223
2 0 12 0 0 8320 0 16 0 0 14 3
366 1345
243 1345
243 1193
1 0 13 0 0 8192 0 16 0 0 13 3
366 1327
333 1327
333 1238
3 1 14 0 0 4224 0 17 14 0 0 3
416 1229
599 1229
599 1219
3 2 13 0 0 12416 0 20 17 0 0 6
559 1000
563 1000
563 1169
291 1169
291 1238
367 1238
3 1 12 0 0 0 0 18 17 0 0 4
223 1193
359 1193
359 1220
367 1220
1 2 11 0 0 0 0 3 18 0 0 4
96 1223
166 1223
166 1202
174 1202
1 1 10 0 0 0 0 4 18 0 0 4
96 1165
166 1165
166 1184
174 1184
3 2 15 0 0 4224 0 21 20 0 0 4
420 1043
505 1043
505 1009
513 1009
3 1 16 0 0 4224 0 22 20 0 0 4
419 969
505 969
505 991
513 991
2 0 17 0 0 4224 0 21 0 0 27 3
375 1052
145 1052
145 843
1 0 18 0 0 4224 0 21 0 0 26 3
375 1034
176 1034
176 895
1 0 19 0 0 8192 0 22 0 0 24 3
374 960
323 960
323 880
2 0 20 0 0 4096 0 22 0 0 25 3
374 978
258 978
258 862
3 1 21 0 0 4224 0 24 23 0 0 3
417 871
659 871
659 864
3 2 19 0 0 12416 0 26 24 0 0 6
588 700
592 700
592 807
295 807
295 880
368 880
3 1 20 0 0 4224 0 25 24 0 0 2
249 862
368 862
1 2 18 0 0 0 0 5 25 0 0 4
137 895
192 895
192 871
200 871
1 1 17 0 0 0 0 6 25 0 0 4
137 843
192 843
192 853
200 853
3 2 22 0 0 4224 0 27 26 0 0 4
452 742
534 742
534 709
542 709
3 1 23 0 0 4224 0 28 26 0 0 4
451 664
534 664
534 691
542 691
0 2 24 0 0 8320 0 0 27 36 0 3
163 575
163 751
407 751
0 1 25 0 0 4224 0 0 27 37 0 3
184 506
184 733
407 733
2 0 26 0 0 8192 0 28 0 0 38 3
406 673
341 673
341 559
1 0 27 0 0 8192 0 28 0 0 35 3
406 655
355 655
355 541
3 1 28 0 0 4224 0 30 29 0 0 3
436 550
648 550
648 547
3 1 27 0 0 4224 0 31 30 0 0 2
264 541
387 541
1 2 24 0 0 0 0 7 31 0 0 4
135 575
207 575
207 550
215 550
1 1 25 0 0 0 0 8 31 0 0 4
132 506
207 506
207 532
215 532
3 2 26 0 0 20608 0 34 30 0 0 8
550 305
591 305
591 304
591 304
591 430
324 430
324 559
387 559
3 1 29 0 0 4224 0 37 32 0 0 3
430 191
642 191
642 188
3 2 30 0 0 4224 0 35 34 0 0 4
431 349
496 349
496 314
504 314
3 1 31 0 0 4224 0 36 34 0 0 4
429 278
496 278
496 296
504 296
0 2 32 0 0 8320 0 0 35 48 0 3
173 181
173 358
386 358
0 1 33 0 0 8320 0 0 35 49 0 3
158 124
158 340
386 340
0 2 2 0 0 4096 0 0 36 46 0 3
305 200
305 287
384 287
0 1 34 0 0 4224 0 0 36 47 0 3
350 179
350 269
384 269
1 2 2 0 0 8320 0 33 37 0 0 3
67 259
67 200
381 200
3 1 34 0 0 0 0 38 37 0 0 4
274 143
350 143
350 182
381 182
1 2 32 0 0 0 0 9 38 0 0 4
134 181
217 181
217 152
225 152
1 1 33 0 0 0 0 10 38 0 0 4
133 124
217 124
217 134
225 134
3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
593 162 622 186
603 170 611 186
1 S
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
587 289 640 313
597 297 629 313
4 Cout
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
83 193 128 217
93 201 117 217
3 Cin
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
