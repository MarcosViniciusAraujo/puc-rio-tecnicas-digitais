CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
260 620 30 90 10
176 80 1278 651
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.440191 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
43
8 2-In OR~
219 724 1003 0 1 22
0 0
0
0 0 608 180
6 74LS32
-21 -24 21 -16
4 U16A
-2 -25 26 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
5130 0 0
2
44899.5 0
0
5 4082~
219 1120 675 0 1 22
0 0
0
0 0 608 270
4 4082
-7 -24 21 -16
4 U15A
20 -4 48 4
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 4 0
1 U
391 0 0
2
44899.5 0
0
13 Logic Switch~
5 57 1011 0 1 11
0 14
0
0 0 21344 0
2 0V
-6 -16 8 -8
4 INIC
-13 -26 15 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.90056e-315 0
0
13 Logic Switch~
5 148 1071 0 1 11
0 18
0
0 0 21344 0
2 0V
-6 -16 8 -8
5 CLOCK
-16 -26 19 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
5.90056e-315 0
0
13 Logic Switch~
5 531 849 0 1 11
0 25
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
5.90056e-315 0
0
9 Inverter~
13 557 1081 0 2 22
0 3 4
0
0 0 608 0
6 74LS04
-21 -19 21 -11
4 U13D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 2 0
1 U
5572 0 0
2
5.90056e-315 0
0
5 4013~
219 627 1102 0 6 22
0 3 3 4 79 80 5
0
0 0 4704 0
4 4013
10 -60 38 -52
4 U14A
23 -61 51 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 3 0
1 U
8901 0 0
2
5.90056e-315 0
0
14 Logic Display~
6 664 1028 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7361 0 0
2
5.90056e-315 0
0
9 Inverter~
13 276 1011 0 2 22
0 14 6
0
0 0 608 0
6 74LS04
-21 -19 21 -11
4 U13C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 2 0
1 U
4747 0 0
2
5.90056e-315 0
0
12 Hex Display~
7 641 872 0 16 19
10 10 9 8 7 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
972 0 0
2
5.90056e-315 0
0
7 Ground~
168 1313 607 0 1 3
0 2
0
0 0 53344 0
0
5 GND11
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3472 0 0
2
5.90056e-315 0
0
2 +V
167 1453 593 0 1 3
0 11
0
0 0 54240 0
2 5V
-7 -22 7 -14
2 V6
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9998 0 0
2
5.90056e-315 0
0
7 Ground~
168 1140 594 0 1 3
0 2
0
0 0 53344 0
0
5 GND10
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3536 0 0
2
5.90056e-315 0
0
7 Ground~
168 1043 637 0 1 3
0 2
0
0 0 53344 0
0
4 GND9
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4597 0 0
2
5.90056e-315 0
0
9 Inverter~
13 923 1133 0 2 22
0 13 12
0
0 0 608 0
6 74LS04
-21 -19 21 -11
4 U13B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
3835 0 0
2
5.90056e-315 0
0
7 Ground~
168 456 711 0 1 3
0 2
0
0 0 53344 0
0
4 GND8
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3670 0 0
2
5.90056e-315 0
0
7 Ground~
168 434 358 0 1 3
0 2
0
0 0 53344 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5616 0 0
2
5.90056e-315 0
0
7 Ground~
168 331 1193 0 1 3
0 2
0
0 0 53344 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9323 0 0
2
5.90056e-315 0
0
7 Ground~
168 796 713 0 1 3
0 2
0
0 0 53344 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
317 0 0
2
5.90056e-315 0
0
7 Ground~
168 790 512 0 1 3
0 2
0
0 0 53344 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3108 0 0
2
5.90056e-315 0
0
7 Ground~
168 284 1106 0 1 3
0 2
0
0 0 53344 180
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4299 0 0
2
5.90056e-315 0
0
2 +V
167 307 1100 0 1 3
0 11
0
0 0 54240 0
2 5V
-7 -22 7 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9672 0 0
2
5.90056e-315 0
0
9 Inverter~
13 370 1052 0 2 22
0 20 19
0
0 0 608 180
6 74LS04
-21 -19 21 -11
4 U13A
-8 -20 20 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
7876 0 0
2
5.90056e-315 0
0
7 Ground~
168 489 1179 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6369 0 0
2
5.90056e-315 0
0
7 74LS191
135 380 1122 0 14 29
0 3 18 19 2 2 2 2 2 81
82 83 20 21 22
0
0 0 4832 0
6 74F191
-21 -51 21 -43
3 U12
-11 -52 10 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 14 11 5 9 10 1 15 13
12 7 6 2 3 4 14 11 5 9
10 1 15 13 12 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
9172 0 0
2
5.90056e-315 0
0
4 4555
219 533 1162 0 7 32
0 21 22 2 17 16 13 15
0
0 0 4832 0
4 4555
-14 -60 14 -52
4 U11A
-14 -61 14 -53
0
15 DVDD=16;DGND=8;
65 %D [%16bi %8bi %1i %2i %3i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 3 2 1 4 5 6 7 3 2
1 4 5 6 7 13 14 15 12 11
10 9 0 0 0 0 0 0 0 0
0 19 0
65 0 0 0 2 1 1 0
1 U
7100 0 0
2
5.90056e-315 0
0
2 +V
167 463 903 0 1 3
0 26
0
0 0 54240 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3820 0 0
2
5.90056e-315 0
0
7 74LS174
130 1393 586 0 14 29
0 16 2 2 27 28 29 30 11 84
85 27 28 29 30
0
0 0 4832 692
7 74LS174
-24 -51 25 -43
3 U10
-11 -53 10 -45
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 9 14 13 11 6 4 3 1 15
12 10 7 5 2 9 14 13 11 6
4 3 1 15 12 10 7 5 2 0
65 0 0 512 1 0 0 0
1 U
7678 0 0
2
5.90056e-315 0
0
7 74LS245
64 1189 543 0 18 37
0 86 87 88 89 31 32 33 34 90
91 92 93 27 28 29 30 2 12
0
0 0 4832 692
7 74LS245
-24 -60 25 -52
2 U9
-7 -62 7 -54
0
16 DVCC=20;DGND=10;
192 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i]
+ [%20bi %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP14
37

0 9 8 7 6 5 4 3 2 11
12 13 14 15 16 17 18 19 1 9
8 7 6 5 4 3 2 11 12 13
14 15 16 17 18 19 1 0
65 0 0 512 1 0 0 0
1 U
961 0 0
2
5.90056e-315 0
0
7 Ground~
168 994 633 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3178 0 0
2
5.90056e-315 0
0
6 1K RAM
79 1031 552 0 20 41
0 2 2 35 36 37 38 39 40 41
42 94 95 96 97 31 32 33 34 2
12
0
0 0 4832 692
5 RAM1K
-17 -19 18 -11
2 U8
-7 -71 7 -63
0
16 DVCC=22;DGND=11;
214 %D [%22bi %11bi  %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i %19i %20i]
+ [%22bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o  %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o] %M
0
12 type:digital
5 DIP22
41

0 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 0
65 0 0 512 1 0 0 0
1 U
3409 0 0
2
5.90056e-315 0
0
7 74LS157
122 835 646 0 14 29
0 13 46 54 45 53 44 52 43 51
2 38 37 36 35
0
0 0 4832 0
6 74F157
-21 -60 21 -52
2 U7
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
3951 0 0
2
5.90056e-315 0
0
7 74LS157
122 837 437 0 14 29
0 13 50 58 49 57 48 56 47 55
2 42 41 40 39
0
0 0 4832 0
6 74F157
-21 -60 21 -52
2 U6
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
8885 0 0
2
5.90056e-315 0
0
7 74LS191
135 547 761 0 14 29
0 2 23 6 2 63 64 65 66 98
99 43 44 45 46
0
0 0 4832 0
6 74F191
-21 -51 21 -43
2 U4
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 14 11 5 9 10 1 15 13
12 7 6 2 3 4 14 11 5 9
10 1 15 13 12 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
3780 0 0
2
5.90056e-315 5.26354e-315
0
7 74LS191
135 553 645 0 14 29
0 2 15 6 2 67 68 69 70 23
100 47 48 49 50
0
0 0 4832 0
6 74F191
-21 -51 21 -43
2 U3
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 14 11 5 9 10 1 15 13
12 7 6 2 3 4 14 11 5 9
10 1 15 13 12 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
9265 0 0
2
5.90056e-315 0
0
7 74LS191
135 549 432 0 14 29
0 2 24 6 2 71 72 73 74 101
102 51 52 53 54
0
0 0 4832 0
6 74F191
-21 -51 21 -43
2 U2
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 14 11 5 9 10 1 15 13
12 7 6 2 3 4 14 11 5 9
10 1 15 13 12 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
9442 0 0
2
5.90056e-315 5.26354e-315
0
7 74LS191
135 546 278 0 14 29
0 2 15 6 2 75 76 77 78 24
103 55 56 57 58
0
0 0 4832 0
6 74F191
-21 -51 21 -43
2 U1
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 14 11 5 9 10 1 15 13
12 7 6 2 3 4 14 11 5 9
10 1 15 13 12 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
9424 0 0
2
5.90056e-315 0
0
7 74LS191
135 539 920 0 14 29
0 25 15 6 26 59 60 61 62 104
3 7 8 9 10
0
0 0 4832 0
6 74F191
-21 -51 21 -43
2 U5
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 14 11 5 9 10 1 15 13
12 7 6 2 3 4 14 11 5 9
10 1 15 13 12 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
9968 0 0
2
5.90056e-315 0
0
8 Hex Key~
166 99 822 0 11 12
0 62 61 60 59 0 0 0 0 0
2 50
0
0 0 4640 0
0
2 NP
-7 -34 7 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
9281 0 0
2
5.90056e-315 0
0
8 Hex Key~
166 101 679 0 11 12
0 66 65 64 63 0 0 0 0 0
0 48
0
0 0 4640 0
0
4 EDF2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
8464 0 0
2
5.90056e-315 0
0
8 Hex Key~
166 101 560 0 11 12
0 70 69 68 67 0 0 0 0 0
10 65
0
0 0 4640 0
0
4 EDF1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
7168 0 0
2
5.90056e-315 0
0
8 Hex Key~
166 102 323 0 11 12
0 74 73 72 71 0 0 0 0 0
0 48
0
0 0 4640 0
0
4 EDI2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3171 0 0
2
5.90056e-315 0
0
8 Hex Key~
166 100 193 0 11 12
0 78 77 76 75 0 0 0 0 0
0 48
0
0 0 4640 0
0
4 EDI1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
4139 0 0
2
5.90056e-315 0
0
164
5 1 0 0 0 0 0 2 1 0 0 3
1118 698
1118 1012
743 1012
3 0 0 0 0 0 0 1 0 0 3 4
697 1003
624 1003
624 1026
619 1026
1 1 0 0 0 12432 0 7 25 0 0 5
627 1045
619 1045
619 1025
342 1025
342 1095
1 0 0 0 0 0 0 2 0 0 77 4
1131 653
1131 606
1126 606
1126 526
2 0 0 0 0 0 0 2 0 0 78 4
1122 653
1122 522
1123 522
1123 517
3 0 0 0 0 0 0 2 0 0 79 2
1113 653
1113 508
4 0 0 0 0 0 0 2 0 0 80 2
1104 653
1104 499
0 0 3 0 0 4100 0 0 0 0 0 3
619 1025
619 1045
627 1045
2 3 4 0 0 4224 0 6 7 0 0 4
578 1081
595 1081
595 1084
603 1084
0 1 3 0 0 4096 0 0 6 3 0 3
530 1025
530 1081
542 1081
6 1 5 0 0 8320 0 7 8 0 0 3
651 1066
664 1066
664 1046
0 2 3 0 0 0 0 0 7 3 0 3
599 1025
599 1066
603 1066
2 3 6 0 0 4096 0 9 38 0 0 4
297 1011
421 1011
421 911
501 911
11 4 7 0 0 4224 0 38 10 0 0 3
571 929
632 929
632 896
12 3 8 0 0 4224 0 38 10 0 0 3
571 938
638 938
638 896
13 2 9 0 0 4224 0 38 10 0 0 3
571 947
644 947
644 896
14 1 10 0 0 4224 0 38 10 0 0 3
571 956
650 956
650 896
2 0 2 0 0 4096 0 28 0 0 19 3
1361 596
1333 596
1333 587
3 1 2 0 0 4096 0 28 11 0 0 3
1361 587
1313 587
1313 601
8 1 11 0 0 4224 0 28 12 0 0 3
1431 605
1453 605
1453 602
18 0 12 0 0 12288 0 29 0 0 24 4
1221 571
1225 571
1225 718
1085 718
17 1 2 0 0 0 0 29 13 0 0 3
1151 571
1140 571
1140 588
19 1 2 0 0 0 0 31 14 0 0 5
1069 580
1073 580
1073 623
1043 623
1043 631
2 20 12 0 0 8320 0 15 31 0 0 4
944 1133
1085 1133
1085 571
1069 571
0 1 13 0 0 4096 0 0 15 50 0 2
757 1133
908 1133
10 2 3 0 0 12432 0 38 1 0 0 4
571 920
765 920
765 994
743 994
0 3 6 0 0 4096 0 0 37 28 0 3
424 424
424 269
508 269
0 3 6 0 0 4224 0 0 36 29 0 3
424 636
424 423
511 423
0 3 6 0 0 0 0 0 35 30 0 3
421 753
421 636
515 636
0 3 6 0 0 0 0 0 34 13 0 3
421 912
421 752
509 752
1 1 14 0 0 4224 0 3 9 0 0 2
69 1011
261 1011
1 0 2 0 0 0 0 36 0 0 38 4
511 405
483 405
483 406
478 406
1 0 2 0 0 0 0 37 0 0 39 4
508 251
503 251
503 278
500 278
1 0 2 0 0 0 0 34 0 0 36 2
509 734
470 734
1 0 2 0 0 0 0 35 0 0 37 3
515 618
467 618
467 645
4 0 2 0 0 8192 0 34 0 0 37 4
515 761
470 761
470 689
456 689
4 1 2 0 0 0 0 35 16 0 0 3
521 645
456 645
456 705
0 4 2 0 0 0 0 0 36 39 0 3
478 366
478 432
517 432
1 4 2 0 0 28800 0 17 37 0 0 9
434 352
434 344
447 344
447 362
457 362
457 366
500 366
500 278
514 278
0 2 15 0 0 4224 0 0 37 41 0 3
492 627
492 260
514 260
0 2 15 0 0 0 0 0 35 46 0 3
492 903
492 627
521 627
8 0 2 0 0 0 0 25 0 0 45 2
348 1158
331 1158
7 0 2 0 0 0 0 25 0 0 45 2
348 1149
331 1149
6 0 2 0 0 0 0 25 0 0 45 2
348 1140
331 1140
5 1 2 0 0 0 0 25 18 0 0 3
348 1131
331 1131
331 1187
7 2 15 0 0 0 0 26 38 0 0 6
565 1135
586 1135
586 1003
492 1003
492 902
507 902
10 1 2 0 0 0 0 32 19 0 0 5
797 691
788 691
788 699
796 699
796 707
10 1 2 0 0 0 0 33 20 0 0 3
799 482
790 482
790 506
0 1 13 0 0 4096 0 0 33 50 0 3
757 612
757 401
805 401
6 1 13 0 0 8320 0 26 32 0 0 4
565 1144
757 1144
757 610
803 610
1 5 16 0 0 12416 0 28 26 0 0 4
1361 605
1336 605
1336 1153
565 1153
4 0 17 0 0 4224 0 26 0 0 0 3
565 1162
602 1162
602 1161
1 2 18 0 0 4224 0 4 25 0 0 4
160 1071
329 1071
329 1104
348 1104
1 4 2 0 0 0 0 21 25 0 0 3
284 1114
284 1122
348 1122
2 3 19 0 0 8320 0 23 25 0 0 4
355 1052
334 1052
334 1113
342 1113
12 1 20 0 0 12416 0 25 23 0 0 5
412 1140
412 1138
422 1138
422 1052
391 1052
13 1 21 0 0 4224 0 25 26 0 0 4
412 1149
482 1149
482 1135
501 1135
14 2 22 0 0 4224 0 25 26 0 0 4
412 1158
488 1158
488 1144
501 1144
3 1 2 0 0 0 0 26 24 0 0 3
495 1162
489 1162
489 1173
9 2 23 0 0 12416 0 35 34 0 0 6
591 636
595 636
595 714
501 714
501 743
515 743
9 2 24 0 0 8320 0 37 36 0 0 6
584 269
591 269
591 385
503 385
503 414
517 414
1 1 25 0 0 8320 0 38 5 0 0 4
501 893
501 858
543 858
543 849
1 4 26 0 0 8320 0 27 38 0 0 3
463 912
463 920
507 920
11 3 27 0 0 12416 0 28 0 0 76 4
1425 578
1490 578
1490 446
1284 446
12 2 28 0 0 12416 0 28 0 0 76 4
1425 569
1475 569
1475 461
1284 461
13 1 29 0 0 12416 0 28 0 0 76 4
1425 560
1458 560
1458 479
1284 479
14 0 30 0 0 12416 0 28 0 0 76 4
1425 551
1438 551
1438 492
1284 492
4 3 27 0 0 0 0 28 0 0 76 2
1361 578
1284 578
5 2 28 0 0 0 0 28 0 0 76 2
1361 569
1284 569
6 1 29 0 0 0 0 28 0 0 76 2
1361 560
1284 560
7 0 30 0 0 0 0 28 0 0 76 2
1361 551
1284 551
13 3 27 0 0 0 0 29 0 0 76 2
1221 526
1284 526
14 2 28 0 0 0 0 29 0 0 76 2
1221 517
1284 517
15 1 29 0 0 0 0 29 0 0 76 2
1221 508
1284 508
16 0 30 0 0 0 0 29 0 0 76 2
1221 499
1284 499
-150640 0 1 0 0 4128 0 0 0 0 0 2
1284 371
1284 704
15 5 31 0 0 4224 0 31 29 0 0 2
1063 526
1157 526
16 6 32 0 0 4224 0 31 29 0 0 2
1063 517
1157 517
17 7 33 0 0 4224 0 31 29 0 0 2
1063 508
1157 508
18 8 34 0 0 4224 0 31 29 0 0 2
1063 499
1157 499
0 1 2 0 0 0 0 0 30 83 0 3
991 580
994 580
994 627
14 3 35 0 0 8320 0 32 31 0 0 4
867 682
978 682
978 562
999 562
2 1 2 0 0 0 0 31 31 0 0 4
999 571
983 571
983 580
999 580
13 4 36 0 0 8320 0 32 31 0 0 4
867 664
969 664
969 553
999 553
12 5 37 0 0 8320 0 32 31 0 0 4
867 646
955 646
955 544
999 544
11 6 38 0 0 8320 0 32 31 0 0 4
867 628
943 628
943 535
999 535
14 7 39 0 0 4224 0 33 31 0 0 4
869 473
934 473
934 526
999 526
13 8 40 0 0 4224 0 33 31 0 0 4
869 455
952 455
952 517
999 517
12 9 41 0 0 4224 0 33 31 0 0 4
869 437
965 437
965 508
999 508
11 10 42 0 0 4224 0 33 31 0 0 4
869 419
977 419
977 499
999 499
8 -154809 43 0 0 12288 0 32 0 0 123 4
803 673
782 673
782 732
711 732
6 -154810 44 0 0 8192 0 32 0 0 123 4
803 655
769 655
769 719
711 719
4 -154811 45 0 0 4096 0 32 0 0 123 2
803 637
711 637
2 -154812 46 0 0 4096 0 32 0 0 123 2
803 619
711 619
8 -154813 47 0 0 4096 0 33 0 0 123 2
805 464
711 464
6 -154814 48 0 0 4096 0 33 0 0 123 2
805 446
711 446
4 -154815 49 0 0 4096 0 33 0 0 123 2
805 428
711 428
2 -154816 50 0 0 4096 0 33 0 0 123 2
805 410
711 410
9 -154489 51 0 0 4096 0 32 0 0 123 4
803 682
748 682
748 714
711 714
7 -154490 52 0 0 4096 0 32 0 0 123 4
803 664
729 664
729 697
711 697
5 -154491 53 0 0 4096 0 32 0 0 123 2
803 646
711 646
3 -154492 54 0 0 4096 0 32 0 0 123 2
803 628
711 628
9 -154493 55 0 0 4096 0 33 0 0 123 2
805 473
711 473
7 -154494 56 0 0 4096 0 33 0 0 123 2
805 455
711 455
5 -154495 57 0 0 4096 0 33 0 0 123 2
805 437
711 437
3 -154496 58 0 0 4096 0 33 0 0 123 2
805 419
711 419
11 -154809 43 0 0 4224 0 34 0 0 123 2
579 770
711 770
12 -154810 44 0 0 4224 0 34 0 0 123 2
579 779
711 779
13 -154811 45 0 0 4224 0 34 0 0 123 2
579 788
711 788
14 -154812 46 0 0 4224 0 34 0 0 123 2
579 797
711 797
11 -154813 47 0 0 4224 0 35 0 0 123 2
585 654
711 654
12 -154814 48 0 0 4224 0 35 0 0 123 2
585 663
711 663
13 -154815 49 0 0 4224 0 35 0 0 123 2
585 672
711 672
14 -154816 50 0 0 4224 0 35 0 0 123 2
585 681
711 681
11 -154489 51 0 0 4224 0 36 0 0 123 2
581 441
711 441
12 -154490 52 0 0 4224 0 36 0 0 123 2
581 450
711 450
13 -154491 53 0 0 4224 0 36 0 0 123 2
581 459
711 459
14 -154492 54 0 0 4224 0 36 0 0 123 2
581 468
711 468
11 -154493 55 0 0 4224 0 37 0 0 123 2
578 287
711 287
12 -154494 56 0 0 4224 0 37 0 0 123 2
578 296
711 296
13 -154495 57 0 0 4224 0 37 0 0 123 2
578 305
711 305
14 -154496 58 0 0 4224 0 37 0 0 123 2
578 314
711 314
-865999395 0 1 0 0 4128 0 0 0 0 0 2
711 152
711 968
5 -58172 59 0 0 4096 0 38 0 0 164 2
507 929
335 929
6 -58173 60 0 0 4096 0 38 0 0 164 2
507 938
335 938
7 -58174 61 0 0 4096 0 38 0 0 164 2
507 947
335 947
8 -58175 62 0 0 4096 0 38 0 0 164 2
507 956
335 956
5 -13052985 63 0 0 4096 0 34 0 0 164 2
515 770
335 770
6 -13052986 64 0 0 4096 0 34 0 0 164 2
515 779
335 779
7 -13052987 65 0 0 4096 0 34 0 0 164 2
515 788
335 788
8 -13052988 66 0 0 4096 0 34 0 0 164 2
515 797
335 797
5 -13052989 67 0 0 4096 0 35 0 0 164 2
521 654
335 654
6 -13052990 68 0 0 4096 0 35 0 0 164 2
521 663
335 663
7 -13052991 69 0 0 4096 0 35 0 0 164 2
521 672
335 672
8 -13052992 70 0 0 4096 0 35 0 0 164 2
521 681
335 681
5 -13052793 71 0 0 4096 0 36 0 0 164 2
517 441
335 441
6 -13052794 72 0 0 4096 0 36 0 0 164 2
517 450
335 450
7 -13052795 73 0 0 4096 0 36 0 0 164 2
517 459
335 459
8 -13052796 74 0 0 4096 0 36 0 0 164 2
517 468
335 468
5 -13052797 75 0 0 4096 0 37 0 0 164 2
514 287
335 287
6 -13052798 76 0 0 4096 0 37 0 0 164 2
514 296
335 296
7 -13052799 77 0 0 4096 0 37 0 0 164 2
514 305
335 305
8 -13052800 78 0 0 4096 0 37 0 0 164 2
514 314
335 314
4 -13052985 63 0 0 8320 0 40 0 0 164 3
92 703
92 744
335 744
3 -13052986 64 0 0 8320 0 40 0 0 164 3
98 703
98 733
335 733
2 -13052987 65 0 0 8320 0 40 0 0 164 3
104 703
104 724
335 724
1 -13052988 66 0 0 8320 0 40 0 0 164 3
110 703
110 714
335 714
4 -13052989 67 0 0 8320 0 41 0 0 164 3
92 584
92 629
335 629
3 -13052990 68 0 0 8320 0 41 0 0 164 3
98 584
98 618
335 618
2 -13052991 69 0 0 8320 0 41 0 0 164 3
104 584
104 607
335 607
1 -13052992 70 0 0 8320 0 41 0 0 164 3
110 584
110 597
335 597
4 -13052793 71 0 0 8320 0 42 0 0 164 3
93 347
93 396
335 396
3 -13052794 72 0 0 8320 0 42 0 0 164 3
99 347
99 379
335 379
2 -13052795 73 0 0 8320 0 42 0 0 164 3
105 347
105 367
335 367
1 -13052796 74 0 0 8320 0 42 0 0 164 3
111 347
111 356
335 356
4 -13052797 75 0 0 8320 0 43 0 0 164 3
91 217
91 251
335 251
3 -13052798 76 0 0 8320 0 43 0 0 164 3
97 217
97 241
335 241
2 -13052799 77 0 0 8320 0 43 0 0 164 3
103 217
103 233
335 233
1 -13052800 78 0 0 8320 0 43 0 0 164 3
109 217
109 225
335 225
4 -58172 59 0 0 8320 0 39 0 0 164 3
90 846
90 902
335 902
3 -58173 60 0 0 8320 0 39 0 0 164 3
96 846
96 897
335 897
2 -58174 61 0 0 8320 0 39 0 0 164 3
102 846
102 892
335 892
1 -58175 62 0 0 8320 0 39 0 0 164 3
108 846
108 888
335 888
-902506802 0 1 0 0 4256 0 0 0 0 0 2
335 144
335 963
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
