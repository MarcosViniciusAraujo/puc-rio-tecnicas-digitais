CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 1 100 10
176 80 1278 651
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
15
13 Logic Switch~
5 236 110 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
44828.7 0
0
13 Logic Switch~
5 436 121 0 1 11
0 18
0
0 0 21360 180
2 0V
-7 -16 7 -8
2 V2
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
44828.7 0
0
7 Ground~
168 595 263 0 1 3
0 2
0
0 0 53360 180
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3124 0 0
2
44828.7 0
0
14 Logic Display~
6 833 275 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3421 0 0
2
44828.7 0
0
6 74LS93
109 661 318 0 8 17
0 2 2 5 4 3 27 28 4
0
0 0 4848 0
6 74LS93
-21 -35 21 -27
2 U4
-7 -36 7 -28
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 512 0 0 0 0
1 U
8157 0 0
2
44828.7 0
0
9 2-In AND~
219 535 306 0 3 22
0 7 6 5
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
5572 0 0
2
44828.7 0
0
2 +V
167 548 91 0 1 3
0 8
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
8901 0 0
2
44828.7 0
0
12 Hex Display~
7 721 103 0 16 19
10 13 12 11 10 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
7361 0 0
2
44828.7 0
0
12 Hex Display~
7 767 103 0 16 19
10 17 16 15 14 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
4747 0 0
2
44828.7 0
0
7 Ground~
168 415 179 0 1 3
0 2
0
0 0 53360 90
0
4 GND1
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
972 0 0
2
44828.7 0
0
7 Pulser~
4 348 70 0 10 12
0 29 30 7 31 0 0 5 5 5
8
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
3472 0 0
2
44828.7 0
0
8 Hex Key~
166 142 133 0 11 12
0 22 21 20 19 0 0 0 0 0
11 66
0
0 0 4656 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
9998 0 0
2
44828.7 0
0
8 Hex Key~
166 179 133 0 11 12
0 26 25 24 23 0 0 0 0 0
13 68
0
0 0 4656 512
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
3536 0 0
2
44828.7 0
0
7 74LS164
127 614 178 0 12 25
0 8 9 7 6 10 11 12 13 14
15 16 17
0
0 0 4848 0
6 74F164
-21 -51 21 -43
2 U2
-7 -52 7 -44
0
15 DVCC=14;DGND=7;
96 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 1 2 8 9 13 12 11 10 6
5 4 3 1 2 8 9 13 12 11
10 6 5 4 3 0
65 0 0 0 0 0 0 0
1 U
4597 0 0
2
44828.7 0
0
7 74LS165
97 305 198 0 14 29
0 19 20 21 22 23 24 25 26 18
6 2 7 32 9
0
0 0 4848 0
7 74LS165
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 6 5 4 3 14 13 12 11 10
1 15 2 7 9 6 5 4 3 14
13 12 11 10 1 15 2 7 9 0
65 0 0 512 0 0 0 0
1 U
3835 0 0
2
44828.7 0
0
31
2 0 2 0 0 4096 0 5 0 0 2 3
629 318
629 309
622 309
1 1 2 0 0 4096 0 3 5 0 0 3
595 271
595 309
629 309
5 1 3 0 0 4224 0 5 4 0 0 3
693 309
833 309
833 293
8 4 4 0 0 12416 0 5 5 0 0 6
693 336
697 336
697 351
615 351
615 336
623 336
3 3 5 0 0 4224 0 6 5 0 0 4
556 306
615 306
615 327
623 327
0 2 6 0 0 4096 0 0 6 10 0 3
424 196
424 315
511 315
0 1 7 0 0 4096 0 0 6 11 0 3
481 164
481 297
511 297
1 1 8 0 0 4224 0 7 14 0 0 3
548 100
548 151
582 151
14 2 9 0 0 4224 0 15 14 0 0 4
337 234
568 234
568 160
582 160
0 4 6 0 0 12432 0 0 14 20 0 4
356 141
361 141
361 196
576 196
0 3 7 0 0 4224 0 0 14 23 0 4
382 164
546 164
546 178
582 178
5 4 10 0 0 4224 0 14 8 0 0 3
646 151
712 151
712 127
6 3 11 0 0 4224 0 14 8 0 0 3
646 160
718 160
718 127
7 2 12 0 0 4224 0 14 8 0 0 3
646 169
724 169
724 127
8 1 13 0 0 4224 0 14 8 0 0 3
646 178
730 178
730 127
9 4 14 0 0 4224 0 14 9 0 0 3
646 187
758 187
758 127
10 3 15 0 0 4224 0 14 9 0 0 3
646 196
764 196
764 127
11 2 16 0 0 4224 0 14 9 0 0 3
646 205
770 205
770 127
12 1 17 0 0 4224 0 14 9 0 0 3
646 214
776 214
776 127
1 10 6 0 0 128 0 1 15 0 0 5
236 122
236 125
356 125
356 171
343 171
1 9 18 0 0 4224 0 2 15 0 0 4
422 121
351 121
351 162
337 162
11 1 2 0 0 4224 0 15 10 0 0 2
343 180
408 180
3 12 7 0 0 128 0 11 15 0 0 4
372 61
382 61
382 189
337 189
4 1 19 0 0 8320 0 12 15 0 0 3
133 157
133 171
273 171
3 2 20 0 0 8320 0 12 15 0 0 3
139 157
139 180
273 180
2 3 21 0 0 8320 0 12 15 0 0 3
145 157
145 189
273 189
1 4 22 0 0 8320 0 12 15 0 0 3
151 157
151 198
273 198
4 5 23 0 0 8320 0 13 15 0 0 3
188 157
188 207
273 207
3 6 24 0 0 8320 0 13 15 0 0 3
182 157
182 216
273 216
2 7 25 0 0 8320 0 13 15 0 0 3
176 157
176 225
273 225
1 8 26 0 0 8320 0 13 15 0 0 3
170 157
170 234
273 234
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
