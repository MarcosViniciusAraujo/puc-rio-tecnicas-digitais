CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
190 40 30 120 10
195 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
363 176 476 273
42991634 0
0
6 Title:
5 Name:
0
0
0
20
13 Logic Switch~
5 293 395 0 1 11
0 12
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
44899.9 0
0
13 Logic Switch~
5 243 273 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
391 0 0
2
44899.9 0
0
13 Logic Switch~
5 291 460 0 1 11
0 20
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3124 0 0
2
44899.9 0
0
12 Hex Display~
7 478 174 0 18 19
10 6 5 4 3 0 0 0 0 0
0 1 0 0 1 1 1 0 12
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
3421 0 0
2
44899.9 0
0
9 Inverter~
13 512 461 0 2 22
0 20 7
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
8157 0 0
2
44899.9 0
0
12 Hex Display~
7 598 177 0 18 19
10 11 10 9 8 0 0 0 0 0
0 1 0 0 0 1 1 1 15
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
5572 0 0
2
44899.9 0
0
9 Inverter~
13 318 353 0 2 22
0 12 13
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U1B
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
8901 0 0
2
44899.9 0
0
7 Ground~
168 321 186 0 1 3
0 2
0
0 0 53360 180
0
4 GND8
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7361 0 0
2
44899.9 0
0
7 Ground~
168 297 255 0 1 3
0 2
0
0 0 53360 270
0
4 GND7
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
4747 0 0
2
44899.9 0
0
7 Ground~
168 463 321 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
972 0 0
2
44899.9 0
0
7 Ground~
168 873 165 0 1 3
0 2
0
0 0 53360 180
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3472 0 0
2
44899.9 0
0
7 Ground~
168 888 293 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
9998 0 0
2
44899.9 0
0
2 +V
167 925 241 0 1 3
0 19
0
0 0 54256 270
2 5V
-7 -15 7 -7
2 V1
-7 -25 7 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3536 0 0
2
44899.9 0
0
4 4008
219 846 238 0 14 29
0 2 2 19 19 3 4 5 6 2
18 17 16 15 21
0
0 0 4848 180
4 4008
-14 -60 14 -52
2 U2
-7 -62 7 -54
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 512 0 0 0 0
1 U
4597 0 0
2
44899.9 0
0
7 Ground~
168 630 309 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3835 0 0
2
44899.9 0
0
7 Ground~
168 312 305 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3670 0 0
2
44899.9 0
0
7 Ground~
168 578 321 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5616 0 0
2
44899.9 0
0
7 74LS245
64 675 265 0 18 37
0 22 23 24 25 8 9 10 11 26
27 28 29 15 16 17 18 2 7
0
0 0 4848 692
6 74F245
-21 -60 21 -52
6 BUFFER
-21 -62 21 -54
0
16 DVCC=20;DGND=10;
192 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i]
+ [%20bi %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP14
37

0 9 8 7 6 5 4 3 2 11
12 13 14 15 16 17 18 19 1 9
8 7 6 5 4 3 2 11 12 13
14 15 16 17 18 19 1 0
65 0 0 512 0 0 0 0
1 U
9323 0 0
2
44899.9 0
0
7 74LS191
135 363 253 0 14 29
0 2 14 13 2 2 2 2 2 30
31 3 4 5 6
0
0 0 4848 692
6 74F191
-21 -51 21 -43
7 COUNTER
-24 -52 25 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 14 11 5 9 10 1 15 13
12 7 6 2 3 4 14 11 5 9
10 1 15 13 12 7 6 2 3 0
65 0 0 512 0 0 0 0
1 U
317 0 0
2
44899.9 0
0
6 1K RAM
79 527 274 0 20 41
0 2 2 2 2 2 2 3 4 5
6 32 33 34 35 8 9 10 11 2
7
0
0 0 4848 692
5 RAM1K
-17 -19 18 -11
3 RAM
-10 -71 11 -63
0
16 DVCC=22;DGND=11;
214 %D [%22bi %11bi  %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i %19i %20i]
+ [%22bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o  %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o] %M
0
12 type:digital
5 DIP22
41

0 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 0
65 0 0 512 0 0 0 0
1 U
3108 0 0
2
44899.9 0
0
54
4 0 3 0 0 4096 0 4 0 0 51 2
469 198
469 248
3 0 4 0 0 4096 0 4 0 0 52 2
475 198
475 239
2 0 5 0 0 4096 0 4 0 0 53 2
481 198
481 230
1 0 6 0 0 4096 0 4 0 0 54 2
487 198
487 221
2 20 7 0 0 12416 0 5 20 0 0 5
533 461
533 460
601 460
601 293
565 293
4 0 8 0 0 4096 0 6 0 0 47 2
589 201
589 248
3 0 9 0 0 4096 0 6 0 0 48 2
595 201
595 239
2 0 10 0 0 4096 0 6 0 0 49 2
601 201
601 230
1 0 11 0 0 4096 0 6 0 0 50 2
607 201
607 221
1 1 12 0 0 4224 0 7 1 0 0 3
321 371
321 395
305 395
3 2 13 0 0 8320 0 19 7 0 0 3
325 266
321 266
321 335
2 1 14 0 0 8320 0 19 2 0 0 3
331 275
331 273
255 273
5 0 2 0 0 4096 0 19 0 0 14 3
331 248
321 248
321 239
6 0 2 0 0 0 0 19 0 0 15 3
331 239
321 239
321 230
7 0 2 0 0 8192 0 19 0 0 16 3
331 230
321 230
321 216
8 1 2 0 0 8192 0 19 8 0 0 3
331 221
321 221
321 194
4 1 2 0 0 0 0 19 9 0 0 3
331 257
331 256
304 256
6 0 2 0 0 0 0 20 0 0 19 3
495 257
489 257
489 266
5 0 2 0 0 0 0 20 0 0 20 3
495 266
486 266
486 275
4 0 2 0 0 0 0 20 0 0 21 3
495 275
480 275
480 284
3 0 2 0 0 0 0 20 0 0 22 3
495 284
474 284
474 293
2 0 2 0 0 0 0 20 0 0 23 3
495 293
468 293
468 302
1 1 2 0 0 4224 0 20 10 0 0 3
495 302
463 302
463 315
13 13 15 0 0 4224 0 14 18 0 0 2
814 248
707 248
12 14 16 0 0 4224 0 14 18 0 0 2
814 239
707 239
11 15 17 0 0 4224 0 14 18 0 0 2
814 230
707 230
10 16 18 0 0 4224 0 14 18 0 0 2
814 221
707 221
1 9 2 0 0 0 0 11 14 0 0 4
873 173
873 179
878 179
878 194
1 0 2 0 0 0 0 14 0 0 30 2
878 266
888 266
2 1 2 0 0 0 0 14 12 0 0 3
878 257
888 257
888 287
0 3 19 0 0 8192 0 0 14 32 0 3
893 239
893 248
878 248
1 4 19 0 0 8320 0 13 14 0 0 3
913 240
913 239
878 239
5 -3389 3 0 0 8192 0 14 0 0 46 3
878 230
928 230
928 131
6 -3390 4 0 0 8192 0 14 0 0 46 3
878 221
913 221
913 131
7 -3391 5 0 0 8192 0 14 0 0 46 3
878 212
902 212
902 131
8 -3392 6 0 0 8192 0 14 0 0 46 3
878 203
888 203
888 131
0 18 7 0 0 0 0 0 18 5 0 4
601 460
717 460
717 293
707 293
17 1 2 0 0 0 0 18 15 0 0 3
637 293
630 293
630 303
1 1 20 0 0 4224 0 3 5 0 0 3
303 460
497 460
497 461
1 1 2 0 0 0 0 19 16 0 0 3
325 284
312 284
312 299
19 1 2 0 0 0 0 20 17 0 0 3
565 302
578 302
578 315
0 -3389 3 0 0 4224 0 0 0 51 46 2
448 248
448 131
0 -3390 4 0 0 4224 0 0 0 52 46 2
433 239
433 131
0 -3391 5 0 0 4096 0 0 0 53 46 2
419 230
419 131
0 -3392 6 0 0 4096 0 0 0 54 46 2
406 221
406 131
-145514 0 1 0 0 4256 0 0 0 0 0 2
311 131
1101 131
15 5 8 0 0 4224 0 20 18 0 0 4
559 248
644 248
644 248
643 248
16 6 9 0 0 4224 0 20 18 0 0 4
559 239
644 239
644 239
643 239
17 7 10 0 0 4224 0 20 18 0 0 4
559 230
644 230
644 230
643 230
18 8 11 0 0 4224 0 20 18 0 0 4
559 221
644 221
644 221
643 221
11 7 3 0 0 0 0 19 20 0 0 2
395 248
495 248
12 8 4 0 0 0 0 19 20 0 0 2
395 239
495 239
13 9 5 0 0 4224 0 19 20 0 0 2
395 230
495 230
14 10 6 0 0 4224 0 19 20 0 0 2
395 221
495 221
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
