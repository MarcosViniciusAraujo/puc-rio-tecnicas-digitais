CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
60 140 4 100 10
176 80 1278 651
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
3 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
16
9 Inverter~
13 523 455 0 2 22
0 5 2
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U3A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 5 0
1 U
5130 0 0
2
44828.6 0
0
14 Logic Display~
6 935 371 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
391 0 0
2
44828.6 0
0
9 Inverter~
13 497 459 0 2 22
0 6 4
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U2F
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 4 0
1 U
3124 0 0
2
44828.6 0
0
9 Inverter~
13 506 323 0 2 22
0 5 10
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U2E
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 4 0
1 U
3421 0 0
2
44828.6 0
0
9 Inverter~
13 442 321 0 2 22
0 7 9
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U2D
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 4 0
1 U
8157 0 0
2
44828.6 0
0
9 Inverter~
13 705 495 0 2 22
0 14 13
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 4 0
1 U
5572 0 0
2
44828.6 0
0
5 4082~
219 561 495 0 5 22
0 2 4 7 8 14
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U1B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 3 0
1 U
8901 0 0
2
44828.6 0
0
9 Inverter~
13 718 244 0 2 22
0 15 12
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 4 0
1 U
7361 0 0
2
44828.6 0
0
5 4082~
219 576 244 0 5 22
0 9 6 10 11 15
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U1A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 3 0
1 U
4747 0 0
2
44828.6 0
0
6 74LS74
17 827 426 0 12 25
0 18 19 12 13 20 21 22 23 3
24 25 26
0
0 0 4848 0
6 74LS74
-21 -60 21 -52
2 U7
-7 -61 7 -53
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 3 2 4 1 11 12 10 13 5
6 9 8 3 2 4 1 11 12 10
13 5 6 9 8 0
65 0 0 512 0 0 0 0
1 U
972 0 0
2
44828.6 0
0
5 4073~
219 264 489 0 4 22
0 8 7 5 16
0
0 0 624 180
4 4073
-7 -24 21 -16
3 U4B
-13 -25 8 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 2 0
1 U
3472 0 0
2
5.90048e-315 0
0
12 Hex Display~
7 584 335 0 16 19
10 8 27 28 29 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP3
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 1 0 0 0
4 DISP
9998 0 0
2
5.90048e-315 0
0
6 74LS93
109 355 539 0 8 17
0 16 16 11 30 8 8 8 8
0
0 0 4848 0
6 74LS93
-21 -35 21 -27
2 U6
-7 -36 7 -28
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 512 1 0 0 0
1 U
3536 0 0
2
5.90048e-315 0
0
12 Hex Display~
7 637 337 0 18 19
10 7 6 5 11 0 0 0 0 0
0 1 1 1 0 0 0 0 7
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
4597 0 0
2
5.90048e-315 0
0
6 74LS93
109 355 413 0 8 17
0 16 16 17 7 11 5 6 7
0
0 0 4848 0
6 74LS93
-21 -35 21 -27
2 U5
-7 -36 7 -28
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 0 1 0 0 0
1 U
3835 0 0
2
5.90048e-315 0
0
7 Pulser~
4 170 425 0 10 12
0 31 32 17 33 0 0 5 5 4
8
0
0 0 4656 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3670 0 0
2
5.90048e-315 0
0
36
2 1 2 0 0 8336 0 1 7 0 0 3
526 473
526 482
537 482
9 1 3 0 0 4224 0 10 2 0 0 3
859 399
935 399
935 389
2 2 4 0 0 8320 0 3 7 0 0 3
500 477
500 491
537 491
0 1 5 0 0 4112 0 0 1 31 0 2
526 413
526 437
0 1 6 0 0 4096 0 0 3 24 0 2
500 422
500 441
0 3 7 0 0 4096 0 0 7 32 0 3
473 432
473 500
537 500
0 4 8 0 0 4096 0 0 7 23 0 3
520 557
520 509
537 509
1 0 5 0 0 4096 0 4 0 0 31 2
509 341
509 413
1 0 7 0 0 4096 0 5 0 0 32 2
445 339
445 432
1 2 9 0 0 4224 0 9 5 0 0 3
552 231
445 231
445 303
0 2 6 0 0 4096 0 0 9 24 0 3
478 422
478 240
552 240
3 2 10 0 0 8320 0 9 4 0 0 3
552 249
509 249
509 305
0 4 11 0 0 4096 0 0 9 30 0 3
537 404
537 258
552 258
2 3 12 0 0 8320 0 8 10 0 0 4
739 244
781 244
781 408
789 408
2 4 13 0 0 8320 0 6 10 0 0 4
726 495
781 495
781 417
789 417
5 1 14 0 0 4224 0 7 6 0 0 2
582 495
690 495
5 1 15 0 0 4224 0 9 8 0 0 2
597 244
703 244
0 2 16 0 0 8192 0 0 13 28 0 3
309 530
309 539
323 539
0 1 16 0 0 0 0 0 15 34 0 3
312 413
312 404
323 404
7 0 8 0 0 0 0 13 0 0 23 2
387 548
387 548
6 0 8 0 0 0 0 13 0 0 23 2
387 539
387 539
5 0 8 0 0 0 0 13 0 0 23 2
387 530
387 530
0 1 8 0 0 4224 0 0 12 29 0 3
391 557
593 557
593 359
7 2 6 0 0 4224 0 15 14 0 0 3
387 422
640 422
640 361
0 3 11 0 0 4096 0 0 13 30 0 5
433 404
433 572
309 572
309 548
317 548
0 3 5 0 0 8192 0 0 11 31 0 3
411 413
411 480
282 480
0 2 7 0 0 0 0 0 11 35 0 3
315 454
315 489
282 489
4 1 16 0 0 12416 0 11 13 0 0 4
237 489
235 489
235 530
323 530
8 1 8 0 0 0 0 13 11 0 0 4
387 557
391 557
391 498
282 498
5 4 11 0 0 4224 0 15 14 0 0 3
387 404
628 404
628 361
6 3 5 0 0 4224 0 15 14 0 0 3
387 413
634 413
634 361
0 1 7 0 0 8320 0 0 14 35 0 4
396 431
396 432
646 432
646 361
0 3 17 0 0 0 0 0 15 36 0 2
317 422
317 422
0 2 16 0 0 0 0 0 15 28 0 3
235 489
235 413
323 413
8 4 7 0 0 0 0 15 15 0 0 6
387 431
396 431
396 454
314 454
314 431
317 431
3 3 17 0 0 4224 0 16 15 0 0 4
194 416
309 416
309 422
317 422
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
