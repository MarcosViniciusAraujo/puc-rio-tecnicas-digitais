CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
720 310 3 100 10
176 80 1278 651
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
48 C:\Program Files\CircuitMaker 2000 Trial\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
45
12 Hex Display~
7 1575 703 0 18 19
10 6 5 4 3 0 0 0 0 0
0 1 1 1 1 0 0 1 3
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP3
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
5130 0 0
2
44899.5 0
0
7 Ground~
168 1361 872 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
391 0 0
2
44899.5 0
0
9 Inverter~
13 1115 704 0 2 22
0 11 8
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U7B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 4 0
1 U
3124 0 0
2
44899.5 0
0
5 4082~
219 1185 708 0 5 22
0 12 8 10 9 7
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U10A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 5 0
1 U
3421 0 0
2
44899.5 0
0
7 74LS157
122 1410 796 0 14 29
0 7 2 9 2 10 2 11 2 12
2 6 5 4 3
0
0 0 4848 0
6 74F157
-21 -60 21 -52
2 U9
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 0 0 0 0
1 U
8157 0 0
2
44899.5 0
0
12 Hex Display~
7 1075 636 0 18 19
10 9 10 11 12 0 0 0 0 0
0 1 1 1 1 0 0 1 3
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
5572 0 0
2
44899.5 0
0
2 +V
167 940 835 0 1 3
0 13
0
0 0 54256 180
2 5V
7 -2 21 6
2 V2
7 -12 21 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
8901 0 0
2
44899.5 0
0
7 Ground~
168 917 819 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7361 0 0
2
44899.5 0
0
4 4008
219 983 766 0 14 29
0 14 15 16 17 2 2 2 13 2
9 10 11 12 46
0
0 0 4848 0
4 4008
-14 -60 14 -52
2 U8
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 512 0 0 0 0
1 U
4747 0 0
2
44899.5 0
0
12 Hex Display~
7 823 643 0 18 19
10 17 16 15 14 0 0 0 0 0
0 1 1 0 1 1 0 1 2
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
972 0 0
2
5.90055e-315 0
0
9 Inverter~
13 669 714 0 2 22
0 19 18
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U7A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
3472 0 0
2
5.90055e-315 0
0
7 74LS190
134 732 732 0 14 29
0 47 18 19 48 22 23 24 25 49
50 14 15 16 17
0
0 0 4848 0
6 74F190
-21 -51 21 -43
2 U6
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 14 11 5 9 10 1 15 13
12 7 6 2 3 4 14 11 5 9
10 1 15 13 12 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
9998 0 0
2
5.90055e-315 0
0
6 74LS93
109 276 750 0 8 17
0 27 51 26 25 22 23 24 25
0
0 0 4848 0
6 74LS93
-21 -35 21 -27
2 U5
-7 -36 7 -28
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 512 1 0 0 0
1 U
3536 0 0
2
5.90055e-315 0
0
9 2-In AND~
219 277 691 0 3 22
0 23 22 27
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U3C
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
4597 0 0
2
5.90055e-315 0
0
12 Hex Display~
7 364 687 0 18 19
10 25 24 23 22 0 0 0 0 0
0 1 1 1 0 1 1 1 10
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
2 id
-8 -38 6 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3835 0 0
2
5.90055e-315 0
0
7 Ground~
168 684 78 0 1 3
0 2
0
0 0 53360 180
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3670 0 0
2
5.90055e-315 0
0
7 Ground~
168 201 389 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5616 0 0
2
5.90055e-315 0
0
2 +V
167 433 606 0 1 3
0 30
0
0 0 54256 180
2 5V
7 -2 21 6
2 V4
7 -12 21 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9323 0 0
2
5.90055e-315 5.39306e-315
0
2 +V
167 247 607 0 1 3
0 31
0
0 0 54256 180
2 5V
7 -2 21 6
2 V3
7 -12 21 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
317 0 0
2
5.90055e-315 5.38788e-315
0
12 Hex Display~
7 576 473 0 18 19
10 21 20 32 33 0 0 0 0 0
0 1 1 1 1 0 0 1 3
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 linha
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3108 0 0
2
5.90055e-315 5.36716e-315
0
4 4518
219 484 578 0 20 32
0 34 30 32 21 20 32 33 0 0
0 0 0 0 0 0 0 0 0 0
3
0
0 0 4848 0
4 4518
-14 -60 14 -52
3 U4B
-11 -61 10 -53
0
15 DVDD=16;DGND=8;
65 %D [%16bi %8bi %1i %2i %3i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 19 0
65 0 0 0 2 2 3 0
1 U
4299 0 0
2
5.90055e-315 5.3568e-315
0
12 Hex Display~
7 397 482 0 18 19
10 29 28 36 35 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
6 coluna
-21 -38 21 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
9672 0 0
2
5.90055e-315 5.34643e-315
0
9 2-In AND~
219 322 475 0 3 22
0 29 28 34
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U3B
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
7876 0 0
2
5.90055e-315 5.32571e-315
0
4 4518
219 312 578 0 20 32
0 26 31 34 29 28 36 35 0 0
0 0 0 0 0 0 0 0 0 0
1
0
0 0 4848 0
4 4518
-14 -60 14 -52
3 U4A
-11 -61 10 -53
0
15 DVDD=16;DGND=8;
65 %D [%16bi %8bi %1i %2i %3i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 19 0
65 0 0 0 2 1 3 0
1 U
6369 0 0
2
5.90055e-315 5.30499e-315
0
9 2-In AND~
219 219 551 0 3 22
0 37 19 26
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
9172 0 0
2
5.90055e-315 5.26354e-315
0
7 Pulser~
4 112 551 0 10 12
0 52 53 37 54 0 0 5 5 2
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
7100 0 0
2
5.90055e-315 0
0
7 74LS139
118 201 323 0 14 29
0 28 29 2 55 56 57 58 38 39
40 59 60 61 62
0
0 0 4848 602
7 74LS139
-24 -51 25 -43
2 U2
48 -3 62 5
0
15 DVCC=16;DGND=8;
113 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+[%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 13 14 15 7 6 5
4 9 10 11 12 3 2 1 13 14
15 7 6 5 4 9 10 11 12 0
65 0 0 512 1 0 0 0
1 U
3820 0 0
2
5.90055e-315 0
0
14 NO PushButton~
191 218 175 0 2 5
0 41 40
0
0 0 4720 0
0
3 S12
-10 -20 11 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
7678 0 0
2
5.90055e-315 5.30499e-315
0
14 NO PushButton~
191 295 176 0 2 5
0 41 39
0
0 0 4720 0
0
3 S11
-10 -20 11 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
961 0 0
2
5.90055e-315 5.26354e-315
0
14 NO PushButton~
191 373 175 0 2 5
0 41 38
0
0 0 4720 0
0
3 S10
-10 -20 11 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3178 0 0
2
5.90055e-315 0
0
14 NO PushButton~
191 375 133 0 2 5
0 42 38
0
0 0 4720 0
0
2 S9
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3409 0 0
2
5.90055e-315 5.30499e-315
0
14 NO PushButton~
191 297 134 0 2 5
0 42 39
0
0 0 4720 0
0
2 S8
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3951 0 0
2
5.90055e-315 5.26354e-315
0
14 NO PushButton~
191 220 133 0 2 5
0 42 40
0
0 0 4720 0
0
2 S7
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
8885 0 0
2
5.90055e-315 0
0
14 NO PushButton~
191 220 92 0 2 5
0 43 40
0
0 0 4720 0
0
2 S6
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3780 0 0
2
5.90055e-315 5.30499e-315
0
14 NO PushButton~
191 297 93 0 2 5
0 43 39
0
0 0 4720 0
0
2 S5
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
9265 0 0
2
5.90055e-315 5.26354e-315
0
14 NO PushButton~
191 375 92 0 2 5
0 43 38
0
0 0 4720 0
0
2 S4
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
9442 0 0
2
5.90055e-315 0
0
14 NO PushButton~
191 376 47 0 2 5
0 44 38
0
0 0 4720 0
0
2 S3
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
9424 0 0
2
5.90055e-315 0
0
14 NO PushButton~
191 298 48 0 2 5
0 44 39
0
0 0 4720 0
0
2 S2
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
9968 0 0
2
5.90055e-315 0
0
14 NO PushButton~
191 221 47 0 2 5
0 44 40
0
0 0 4720 0
0
2 S1
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
9281 0 0
2
5.90055e-315 0
0
2 +V
167 51 46 0 1 3
0 45
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8464 0 0
2
5.90055e-315 0
0
7 74LS153
119 635 160 0 14 29
0 63 64 65 66 20 21 41 42 43
44 67 2 68 19
0
0 0 4848 692
7 74LS153
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 4 5 6 2 14 13 12 11
10 1 15 7 9 3 4 5 6 2
14 13 12 11 10 1 15 7 9 0
65 0 0 512 1 0 0 0
1 U
7168 0 0
2
5.90055e-315 0
0
9 Resistor~
219 93 201 0 3 5
0 45 41 1
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 18
82 0 0 0 1 0 0 0
1 R
3171 0 0
2
5.90055e-315 0
0
9 Resistor~
219 91 157 0 3 5
0 45 42 1
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 18
82 0 0 0 1 0 0 0
1 R
4139 0 0
2
5.90055e-315 0
0
9 Resistor~
219 93 117 0 3 5
0 45 43 1
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 62
82 0 0 0 1 0 0 0
1 R
6435 0 0
2
5.90055e-315 0
0
9 Resistor~
219 93 71 0 3 5
0 45 44 1
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 74
82 0 0 0 1 0 0 0
1 R
5283 0 0
2
5.90055e-315 0
0
109
4 14 3 0 0 8320 0 1 5 0 0 3
1566 727
1566 832
1442 832
3 13 4 0 0 8320 0 1 5 0 0 3
1572 727
1572 814
1442 814
2 12 5 0 0 8320 0 1 5 0 0 3
1578 727
1578 796
1442 796
1 11 6 0 0 8320 0 1 5 0 0 3
1584 727
1584 778
1442 778
5 1 7 0 0 4240 0 4 5 0 0 4
1206 708
1364 708
1364 760
1378 760
6 0 2 0 0 4096 0 5 0 0 8 2
1378 805
1363 805
4 0 2 0 0 0 0 5 0 0 8 2
1378 787
1363 787
0 2 2 0 0 4224 0 0 5 9 0 3
1363 823
1363 769
1378 769
8 0 2 0 0 0 0 5 0 0 10 3
1378 823
1361 823
1361 841
10 1 2 0 0 0 0 5 2 0 0 3
1372 841
1361 841
1361 866
2 2 8 0 0 4224 0 3 4 0 0 2
1136 704
1161 704
4 0 9 0 0 4096 0 4 0 0 23 2
1161 722
1084 722
3 0 10 0 0 4096 0 4 0 0 22 2
1161 713
1078 713
0 1 11 0 0 4096 0 0 3 21 0 2
1072 704
1100 704
0 1 12 0 0 4096 0 0 4 20 0 2
1066 695
1161 695
0 9 12 0 0 8320 0 0 5 20 0 3
1066 748
1066 832
1378 832
0 7 11 0 0 8320 0 0 5 21 0 3
1069 757
1069 814
1378 814
0 5 10 0 0 8320 0 0 5 22 0 3
1076 766
1076 796
1378 796
0 3 9 0 0 8320 0 0 5 23 0 3
1083 775
1083 778
1378 778
13 4 12 0 0 128 0 9 6 0 0 3
1015 748
1066 748
1066 660
12 3 11 0 0 128 0 9 6 0 0 3
1015 757
1072 757
1072 660
11 2 10 0 0 128 0 9 6 0 0 3
1015 766
1078 766
1078 660
10 1 9 0 0 128 0 9 6 0 0 3
1015 775
1084 775
1084 660
1 8 13 0 0 4224 0 7 9 0 0 3
940 820
940 793
951 793
0 5 2 0 0 0 0 0 9 26 0 4
917 775
943 775
943 766
951 766
0 6 2 0 0 128 0 0 9 27 0 3
917 802
917 775
951 775
0 7 2 0 0 0 0 0 9 28 0 4
917 802
943 802
943 784
951 784
1 9 2 0 0 0 0 8 9 0 0 3
917 813
917 802
951 802
0 1 14 0 0 8320 0 0 9 33 0 3
813 741
813 730
951 730
0 2 15 0 0 8320 0 0 9 34 0 3
818 750
818 739
951 739
0 3 16 0 0 8320 0 0 9 35 0 3
825 759
825 748
951 748
0 4 17 0 0 8320 0 0 9 36 0 3
832 768
832 757
951 757
11 4 14 0 0 128 0 12 10 0 0 3
764 741
814 741
814 667
12 3 15 0 0 128 0 12 10 0 0 3
764 750
820 750
820 667
13 2 16 0 0 128 0 12 10 0 0 3
764 759
826 759
826 667
14 1 17 0 0 128 0 12 10 0 0 3
764 768
832 768
832 667
2 2 18 0 0 4224 0 11 12 0 0 2
690 714
700 714
0 1 19 0 0 4096 0 0 11 39 0 2
638 714
654 714
0 3 19 0 0 4096 0 0 12 58 0 3
638 639
638 723
694 723
0 5 20 0 0 4224 0 0 41 66 0 3
543 569
543 164
603 164
6 0 21 0 0 8320 0 41 0 0 67 3
603 155
530 155
530 578
0 5 22 0 0 4224 0 0 12 47 0 2
353 741
700 741
0 6 23 0 0 4224 0 0 12 48 0 2
359 750
700 750
0 7 24 0 0 4224 0 0 12 49 0 2
365 759
700 759
0 8 25 0 0 4224 0 0 12 50 0 2
373 768
700 768
0 0 22 0 0 0 0 0 0 51 47 3
335 735
335 741
341 741
5 4 22 0 0 0 0 13 15 0 0 3
308 741
355 741
355 711
6 3 23 0 0 0 0 13 15 0 0 3
308 750
361 750
361 711
7 2 24 0 0 0 0 13 15 0 0 3
308 759
367 759
367 711
8 1 25 0 0 0 0 13 15 0 0 3
308 768
373 768
373 711
2 0 22 0 0 0 0 14 0 0 0 3
295 682
335 682
335 742
1 0 23 0 0 0 0 14 0 0 48 3
295 700
318 700
318 750
0 4 25 0 0 0 0 0 13 50 0 6
319 768
312 768
312 783
230 783
230 768
238 768
0 3 26 0 0 12416 0 0 13 76 0 5
244 551
244 590
225 590
225 759
238 759
3 1 27 0 0 8320 0 14 13 0 0 5
250 691
230 691
230 742
244 742
244 741
12 1 2 0 0 128 0 41 16 0 0 3
673 119
684 119
684 86
3 1 2 0 0 0 0 27 17 0 0 4
203 363
203 375
201 375
201 383
14 2 19 0 0 8320 0 41 25 0 0 6
667 137
677 137
677 639
187 639
187 560
195 560
0 1 28 0 0 12416 0 0 27 74 0 5
355 466
351 466
351 376
221 376
221 357
0 2 29 0 0 12416 0 0 27 75 0 5
349 484
346 484
346 371
212 371
212 357
2 1 30 0 0 8320 0 21 18 0 0 3
446 560
433 560
433 591
2 1 31 0 0 8320 0 24 19 0 0 3
274 560
247 560
247 592
0 3 32 0 0 8320 0 0 21 65 0 5
533 560
533 505
438 505
438 578
452 578
7 4 33 0 0 8320 0 21 20 0 0 3
516 551
567 551
567 497
6 3 32 0 0 0 0 21 20 0 0 3
516 560
573 560
573 497
5 2 20 0 0 0 0 21 20 0 0 3
516 569
579 569
579 497
4 1 21 0 0 0 0 21 20 0 0 3
516 578
585 578
585 497
0 1 34 0 0 4224 0 0 21 73 0 4
266 512
429 512
429 551
452 551
7 4 35 0 0 8320 0 24 22 0 0 3
344 551
388 551
388 506
6 3 36 0 0 8320 0 24 22 0 0 3
344 560
394 560
394 506
2 0 28 0 0 0 0 22 0 0 74 4
400 506
400 568
353 568
353 569
1 0 29 0 0 0 0 22 0 0 75 3
406 506
406 578
347 578
3 3 34 0 0 0 0 23 24 0 0 4
295 475
266 475
266 578
280 578
5 2 28 0 0 0 0 24 23 0 0 4
344 569
355 569
355 466
340 466
4 1 29 0 0 0 0 24 23 0 0 4
344 578
349 578
349 484
340 484
3 1 26 0 0 0 0 25 24 0 0 2
240 551
280 551
1 3 37 0 0 4224 0 25 26 0 0 2
195 542
136 542
0 2 38 0 0 8192 0 0 37 79 0 4
350 100
346 100
346 55
359 55
0 2 38 0 0 0 0 0 36 80 0 4
345 141
350 141
350 100
358 100
0 2 38 0 0 0 0 0 31 81 0 4
348 183
345 183
345 141
358 141
8 2 38 0 0 8320 0 27 30 0 0 5
221 287
221 251
348 251
348 183
356 183
0 2 39 0 0 8192 0 0 38 83 0 4
272 101
268 101
268 56
281 56
0 2 39 0 0 0 0 0 35 84 0 4
263 142
272 142
272 101
280 101
0 2 39 0 0 0 0 0 32 85 0 3
263 184
263 142
280 142
2 9 39 0 0 16512 0 29 27 0 0 5
278 184
263 184
263 232
212 232
212 287
0 2 40 0 0 8192 0 0 39 87 0 4
195 100
191 100
191 55
204 55
0 2 40 0 0 0 0 0 34 88 0 4
190 141
195 141
195 100
203 100
0 2 40 0 0 0 0 0 33 89 0 4
193 183
190 183
190 141
203 141
10 2 40 0 0 12416 0 27 28 0 0 5
203 287
203 263
193 263
193 183
201 183
1 0 41 0 0 8192 0 30 0 0 102 3
390 183
394 183
394 201
1 0 41 0 0 0 0 29 0 0 102 3
312 184
316 184
316 201
1 0 41 0 0 0 0 28 0 0 102 3
235 183
239 183
239 201
1 0 42 0 0 8192 0 31 0 0 103 3
392 141
396 141
396 157
1 0 42 0 0 0 0 32 0 0 103 3
314 142
318 142
318 157
1 0 42 0 0 0 0 33 0 0 103 3
237 141
241 141
241 157
1 0 43 0 0 8192 0 36 0 0 104 3
392 100
396 100
396 117
1 0 43 0 0 0 0 35 0 0 104 3
314 101
318 101
318 117
1 0 43 0 0 0 0 34 0 0 104 3
237 100
241 100
241 117
1 0 44 0 0 8192 0 37 0 0 105 3
393 55
397 55
397 71
1 0 44 0 0 0 0 38 0 0 105 3
315 56
319 56
319 71
1 0 44 0 0 0 0 39 0 0 105 3
238 55
242 55
242 71
2 7 41 0 0 4224 0 42 41 0 0 4
111 201
573 201
573 146
603 146
2 8 42 0 0 4224 0 43 41 0 0 4
109 157
558 157
558 137
603 137
2 9 43 0 0 4224 0 44 41 0 0 4
111 117
582 117
582 128
603 128
2 10 44 0 0 4224 0 45 41 0 0 3
111 71
603 71
603 119
0 1 45 0 0 12416 0 0 42 107 0 5
51 157
51 137
50 137
50 201
75 201
0 1 45 0 0 0 0 0 43 108 0 3
51 117
51 157
73 157
0 1 45 0 0 0 0 0 44 109 0 3
51 71
51 117
75 117
1 1 45 0 0 0 0 40 45 0 0 3
51 55
51 71
75 71
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
