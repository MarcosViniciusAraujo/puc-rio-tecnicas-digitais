CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1278 651
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
31
13 Logic Switch~
5 509 433 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
14 0 28 8
3 V16
10 -10 31 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3465 0 0
2
44809.4 0
0
13 Logic Switch~
5 734 438 0 1 11
0 16
0
0 0 21360 90
2 0V
14 0 28 8
3 V15
10 -10 31 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
8396 0 0
2
44809.3 0
0
13 Logic Switch~
5 679 437 0 1 11
0 15
0
0 0 21360 90
2 0V
14 0 28 8
3 V14
10 -10 31 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3685 0 0
2
44809.3 0
0
13 Logic Switch~
5 544 433 0 1 11
0 9
0
0 0 21360 90
2 0V
14 0 28 8
3 V13
10 -10 31 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
7849 0 0
2
44809.3 0
0
13 Logic Switch~
5 630 435 0 1 11
0 14
0
0 0 21360 90
2 0V
14 0 28 8
3 V12
10 -10 31 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
6343 0 0
2
44809.3 0
0
13 Logic Switch~
5 582 433 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
14 0 28 8
3 V11
10 -10 31 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7376 0 0
2
44809.3 0
0
13 Logic Switch~
5 11 98 0 10 11
0 19 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
3 V10
-10 -31 11 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9156 0 0
2
44809.3 0
0
13 Logic Switch~
5 16 354 0 10 11
0 20 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V9
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5776 0 0
2
44809.3 0
0
13 Logic Switch~
5 204 359 0 10 11
0 25 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V8
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7207 0 0
2
44809.3 0
0
13 Logic Switch~
5 150 359 0 10 11
0 24 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V7
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4459 0 0
2
44809.3 0
0
13 Logic Switch~
5 93 359 0 10 11
0 23 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V6
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3760 0 0
2
44809.3 0
0
13 Logic Switch~
5 49 354 0 10 11
0 22 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V5
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
754 0 0
2
44809.3 0
0
13 Logic Switch~
5 53 111 0 10 11
0 26 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9767 0 0
2
44809.3 0
0
13 Logic Switch~
5 100 111 0 1 11
0 27
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
7978 0 0
2
44809.3 0
0
13 Logic Switch~
5 135 114 0 10 11
0 28 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3142 0 0
2
44809.3 0
0
13 Logic Switch~
5 171 113 0 10 11
0 29 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3284 0 0
2
44809.3 0
0
14 Logic Display~
6 389 44 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
659 0 0
2
44809.4 0
0
14 Logic Display~
6 421 48 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3800 0 0
2
44809.3 0
0
14 Logic Display~
6 449 50 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6792 0 0
2
44809.3 0
0
14 Logic Display~
6 475 52 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3701 0 0
2
44809.3 0
0
14 Logic Display~
6 500 53 0 1 2
10 17
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6316 0 0
2
44809.3 0
0
14 Logic Display~
6 526 59 0 1 2
10 18
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8734 0 0
2
44809.3 0
0
7 Ground~
168 851 135 0 1 3
0 2
0
0 0 53360 90
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7988 0 0
2
44809.3 0
0
7 Ground~
168 1013 344 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3217 0 0
2
44809.3 0
0
14 Logic Display~
6 869 411 0 1 2
10 8
0
0 0 53856 180
6 100MEG
3 -16 45 -8
2 L6
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3965 0 0
2
44809.3 0
0
6 74LS85
106 904 265 0 14 29
0 2 2 3 7 2 2 4 9 12
11 10 30 31 8
0
0 0 5104 512
5 74F85
-18 -52 17 -44
2 U4
-7 -62 7 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 0 0 0 0
1 U
8239 0 0
2
44809.3 0
0
6 74LS85
106 739 267 0 14 29
0 5 6 17 18 13 14 15 16 2
2 2 12 11 10
0
0 0 5104 0
5 74F85
-18 -52 17 -44
2 U3
-7 -62 7 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 0 0 0 0 0
1 U
828 0 0
2
44809.3 0
0
7 Ground~
168 211 481 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
6187 0 0
2
44809.3 0
0
4 4008
219 353 422 0 14 29
0 2 2 2 20 2 2 2 19 21
7 3 32 33 34
0
0 0 4848 0
4 4008
-14 -60 14 -52
2 U2
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 512 0 0 0 0
1 U
7107 0 0
2
44809.3 0
0
7 Ground~
168 250 274 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
6433 0 0
2
44809.3 0
0
4 4008
219 269 205 0 14 29
0 26 27 28 29 22 23 24 25 2
18 17 6 5 21
0
0 0 4848 0
4 4008
-14 -60 14 -52
2 U1
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 0 0 0 0 0
1 U
8559 0 0
2
44809.3 0
0
49
0 3 3 0 0 4240 0 0 26 2 0 4
389 122
991 122
991 256
936 256
11 1 3 0 0 128 0 29 17 0 0 3
385 422
389 422
389 62
1 7 4 0 0 8320 0 1 26 0 0 5
510 420
510 328
949 328
949 292
936 292
0 1 5 0 0 8192 0 0 19 40 0 3
468 129
449 129
449 68
0 1 6 0 0 8192 0 0 20 39 0 5
513 102
492 102
492 76
475 76
475 70
0 4 7 0 0 4224 0 0 26 7 0 4
413 154
949 154
949 265
936 265
10 1 7 0 0 0 0 29 18 0 0 5
385 431
413 431
413 115
421 115
421 66
1 0 2 0 0 4096 0 29 0 0 32 3
321 386
224 386
224 440
0 11 2 0 0 0 0 0 27 10 0 3
779 249
779 258
771 258
0 10 2 0 0 0 0 0 27 11 0 3
779 240
779 249
771 249
1 9 2 0 0 8192 0 23 27 0 0 4
844 136
779 136
779 240
771 240
0 1 2 0 0 0 0 0 26 15 0 4
1013 293
1014 293
1014 238
936 238
0 2 2 0 0 0 0 0 26 15 0 3
1007 292
1007 247
936 247
0 5 2 0 0 0 0 0 26 15 0 3
975 292
975 274
936 274
6 1 2 0 0 0 0 26 24 0 0 5
936 283
954 283
954 292
1013 292
1013 338
14 1 8 0 0 8320 0 26 25 0 0 3
872 301
869 301
869 397
1 8 9 0 0 8320 0 4 26 0 0 5
545 420
545 323
944 323
944 301
936 301
14 11 10 0 0 4224 0 27 26 0 0 4
771 303
854 303
854 256
872 256
13 10 11 0 0 4224 0 27 26 0 0 4
771 294
859 294
859 247
872 247
12 9 12 0 0 4224 0 27 26 0 0 4
771 285
864 285
864 238
872 238
1 5 13 0 0 4224 0 6 27 0 0 3
583 420
583 276
707 276
1 6 14 0 0 4224 0 5 27 0 0 3
631 422
631 285
707 285
1 7 15 0 0 4224 0 3 27 0 0 3
680 424
680 294
707 294
1 8 16 0 0 4224 0 2 27 0 0 5
735 425
735 317
699 317
699 303
707 303
0 1 5 0 0 4224 0 0 27 40 0 4
468 185
684 185
684 240
707 240
0 2 6 0 0 4096 0 0 27 39 0 4
506 195
689 195
689 249
707 249
0 3 17 0 0 4096 0 0 27 38 0 4
536 205
694 205
694 258
707 258
0 4 18 0 0 4096 0 0 27 37 0 4
574 214
699 214
699 267
707 267
2 0 2 0 0 0 0 29 0 0 32 3
321 395
247 395
247 440
3 0 2 0 0 0 0 29 0 0 32 3
321 404
267 404
267 440
5 0 2 0 0 0 0 29 0 0 32 3
321 422
292 422
292 440
0 6 2 0 0 0 0 0 29 33 0 4
211 440
313 440
313 431
321 431
1 7 2 0 0 8320 0 28 29 0 0 3
211 475
211 440
321 440
1 8 19 0 0 20608 0 7 29 0 0 6
11 110
10 110
10 333
-1 333
-1 449
321 449
1 4 20 0 0 16512 0 8 29 0 0 5
17 341
17 338
2 338
2 413
321 413
14 9 21 0 0 8320 0 31 29 0 0 6
301 169
311 169
311 355
259 355
259 458
321 458
1 10 18 0 0 16512 0 22 31 0 0 5
526 77
526 95
574 95
574 214
301 214
1 11 17 0 0 20608 0 21 31 0 0 6
500 71
519 71
519 179
536 179
536 205
301 205
0 12 6 0 0 16512 0 0 31 0 0 5
513 95
513 178
506 178
506 196
301 196
13 0 5 0 0 128 0 31 0 0 0 3
301 187
468 187
468 125
9 1 2 0 0 0 0 31 30 0 0 5
237 241
233 241
233 260
250 260
250 268
1 5 22 0 0 8320 0 12 31 0 0 3
50 341
50 205
237 205
1 6 23 0 0 8320 0 11 31 0 0 3
94 346
94 214
237 214
1 7 24 0 0 4224 0 10 31 0 0 3
151 346
151 223
237 223
1 8 25 0 0 4224 0 9 31 0 0 3
205 346
205 232
237 232
1 1 26 0 0 8320 0 13 31 0 0 3
53 123
53 169
237 169
1 2 27 0 0 8320 0 14 31 0 0 3
100 123
100 178
237 178
1 3 28 0 0 8320 0 15 31 0 0 3
135 126
135 187
237 187
1 4 29 0 0 4224 0 16 31 0 0 3
171 125
171 196
237 196
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
