CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 30 5 100 10
176 80 1278 651
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
16
13 Logic Switch~
5 127 99 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.9005e-315 0
0
5 4082~
219 391 491 0 5 22
0 4 5 6 7 8
0
0 0 608 90
4 4082
-7 -24 21 -16
3 U6A
19 -5 40 3
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 4 0
1 U
391 0 0
2
5.9005e-315 0
0
9 Inverter~
13 184 378 0 2 22
0 9 4
0
0 0 608 270
6 74LS04
-21 -19 21 -11
3 U3C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
3124 0 0
2
5.9005e-315 0
0
9 4-In NOR~
219 286 502 0 5 22
0 4 10 7 11 12
0
0 0 608 90
4 4002
-14 -24 14 -16
3 U5A
29 -2 50 6
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
11 typeDigital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 9 0
65 0 0 0 2 1 3 0
1 U
3421 0 0
2
5.9005e-315 0
0
9 2-In NOR~
219 341 406 0 3 22
0 12 8 13
0
0 0 608 90
6 74LS02
-21 -24 21 -16
3 U4A
31 0 52 8
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
8157 0 0
2
5.9005e-315 0
0
9 Inverter~
13 249 146 0 2 22
0 9 14
0
0 0 608 270
6 74LS04
-21 -19 21 -11
3 U3B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
5572 0 0
2
5.9005e-315 0
0
7 Ground~
168 509 322 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8901 0 0
2
5.9005e-315 0
0
7 Ground~
168 324 149 0 1 3
0 2
0
0 0 53344 180
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7361 0 0
2
5.9005e-315 0
0
7 Ground~
168 329 236 0 1 3
0 2
0
0 0 53344 270
0
4 GND1
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4747 0 0
2
5.9005e-315 0
0
2 +V
167 299 267 0 1 3
0 15
0
0 0 54240 90
2 5V
-7 -15 7 -7
2 V3
-7 -25 7 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
972 0 0
2
5.9005e-315 0
0
12 Hex Display~
7 801 99 0 18 19
10 6 5 16 10 0 0 0 0 0
0 1 1 1 1 1 1 1 8
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3472 0 0
2
5.9005e-315 0
0
12 Hex Display~
7 754 100 0 18 19
10 11 7 18 17 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
9998 0 0
2
5.9005e-315 0
0
9 Inverter~
13 503 229 0 2 22
0 20 19
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U3A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
3536 0 0
2
5.9005e-315 0
0
7 74LS190
134 587 270 0 14 29
0 19 3 13 9 2 2 9 2 21
22 17 18 7 11
0
0 0 4832 0
6 74F190
-21 -51 21 -43
2 U2
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 14 11 5 9 10 1 15 13
12 7 6 2 3 4 14 11 5 9
10 1 15 13 12 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
4597 0 0
2
5.9005e-315 0
0
7 Pulser~
4 143 216 0 10 12
0 23 24 3 25 0 0 5 5 5
8
0
0 0 4640 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3835 0 0
2
5.9005e-315 0
0
7 74LS190
134 410 229 0 14 29
0 2 3 13 9 2 14 15 15 26
20 10 16 5 6
0
0 0 4832 0
6 74F190
-21 -51 21 -43
2 U1
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 14 11 5 9 10 1 15 13
12 7 6 2 3 4 14 11 5 9
10 1 15 13 12 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
3670 0 0
2
5.9005e-315 0
0
37
0 2 3 0 0 8192 0 0 14 27 0 5
368 211
368 285
526 285
526 252
555 252
0 1 4 0 0 8192 0 0 2 7 0 4
278 534
278 550
377 550
377 512
2 0 5 0 0 12416 0 2 0 0 30 4
386 512
386 525
462 525
462 256
3 14 6 0 0 12288 0 2 16 0 0 5
395 512
395 517
456 517
456 265
442 265
0 4 7 0 0 4096 0 0 2 10 0 2
404 539
404 512
5 2 8 0 0 8320 0 2 5 0 0 4
390 467
390 440
356 440
356 425
2 1 4 0 0 4224 0 3 4 0 0 4
187 396
187 534
279 534
279 525
0 1 9 0 0 4096 0 0 3 23 0 2
187 182
187 360
2 0 10 0 0 12288 0 4 0 0 28 4
288 525
288 544
451 544
451 238
3 0 7 0 0 8320 0 4 0 0 34 4
297 525
297 539
642 539
642 297
4 0 11 0 0 8320 0 4 0 0 35 4
306 525
306 534
660 534
660 306
5 1 12 0 0 8320 0 4 5 0 0 4
292 469
292 440
338 440
338 425
0 3 13 0 0 4096 0 0 14 14 0 4
347 320
496 320
496 261
549 261
3 3 13 0 0 4224 0 5 16 0 0 3
347 373
347 220
372 220
5 0 2 0 0 4096 0 14 0 0 18 3
555 279
536 279
536 288
8 1 2 0 0 4096 0 14 7 0 0 4
555 306
555 305
509 305
509 316
7 0 9 0 0 8192 0 14 0 0 24 4
555 297
467 297
467 99
339 99
6 0 2 0 0 0 0 14 0 0 16 5
555 288
536 288
536 306
531 306
531 305
2 6 14 0 0 8320 0 6 16 0 0 3
252 164
252 247
378 247
0 1 9 0 0 0 0 0 6 24 0 2
252 99
252 128
0 7 15 0 0 8192 0 0 16 22 0 3
359 265
359 256
378 256
1 8 15 0 0 4224 0 10 16 0 0 2
310 265
378 265
0 4 9 0 0 8320 0 0 14 24 0 5
173 99
173 182
531 182
531 270
555 270
1 4 9 0 0 0 0 1 16 0 0 4
139 99
340 99
340 229
378 229
1 1 2 0 0 8336 0 8 16 0 0 3
324 157
324 202
372 202
1 5 2 0 0 0 0 9 16 0 0 4
336 237
364 237
364 238
378 238
3 2 3 0 0 8320 0 15 16 0 0 5
167 207
167 210
364 210
364 211
378 211
11 4 10 0 0 12416 0 16 11 0 0 5
442 238
484 238
484 146
792 146
792 123
12 3 16 0 0 12416 0 16 11 0 0 5
442 247
535 247
535 141
798 141
798 123
13 2 5 0 0 0 0 16 11 0 0 5
442 256
540 256
540 136
804 136
804 123
14 1 6 0 0 12416 0 16 11 0 0 5
442 265
545 265
545 131
810 131
810 123
11 4 17 0 0 8320 0 14 12 0 0 3
619 279
745 279
745 124
12 3 18 0 0 8320 0 14 12 0 0 3
619 288
751 288
751 124
2 13 7 0 0 0 0 12 14 0 0 3
757 124
757 297
619 297
1 14 11 0 0 0 0 12 14 0 0 3
763 124
763 306
619 306
2 1 19 0 0 12416 0 13 14 0 0 4
524 229
532 229
532 243
549 243
10 1 20 0 0 4224 0 16 13 0 0 2
442 229
488 229
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
