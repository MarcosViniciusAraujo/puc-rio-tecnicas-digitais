CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 120 10
176 80 1278 651
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
5 4 0.500000 0.181488
344 176 457 273
9437202 256
0
2 

2 

0
0
0
21
13 Logic Switch~
5 419 69 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 E
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
44799.7 0
0
13 Logic Switch~
5 335 67 0 1 11
0 14
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 D
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
44799.7 1
0
13 Logic Switch~
5 247 70 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 C
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
44799.7 2
0
13 Logic Switch~
5 163 70 0 1 11
0 13
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 B
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
44799.7 3
0
13 Logic Switch~
5 76 70 0 1 11
0 17
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 A
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
44799.7 4
0
14 Logic Display~
6 540 54 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5572 0 0
2
5.90044e-315 0
0
5 4071~
219 1350 720 0 3 22
0 5 4 3
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U7A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 7 0
1 U
8901 0 0
2
5.90044e-315 5.26354e-315
0
8 4-In OR~
219 1197 603 0 5 22
0 8 7 6 2 5
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U6A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 6 0
1 U
7361 0 0
2
5.90044e-315 5.30499e-315
0
5 4069~
219 567 918 0 2 22
0 13 12
0
0 0 624 0
4 4069
-7 -24 21 -16
3 U5C
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 3 5 0
1 U
4747 0 0
2
5.90044e-315 5.32571e-315
0
5 4069~
219 567 828 0 2 22
0 14 10
0
0 0 624 0
4 4069
-7 -24 21 -16
3 U5B
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 2 5 0
1 U
972 0 0
2
5.90044e-315 5.34643e-315
0
5 4069~
219 567 783 0 2 22
0 13 15
0
0 0 624 0
4 4069
-7 -24 21 -16
3 U5A
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 1 5 0
1 U
3472 0 0
2
5.90044e-315 5.3568e-315
0
5 4049~
219 564 744 0 2 22
0 17 16
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3F
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 3 0
1 U
9998 0 0
2
44799.7 5
0
5 4082~
219 768 756 0 5 22
0 16 15 11 10 2
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U4B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 4 0
1 U
3536 0 0
2
44799.7 6
0
5 4082~
219 768 969 0 5 22
0 12 11 10 9 4
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U4A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 4 0
1 U
4597 0 0
2
44799.7 7
0
5 4049~
219 564 432 0 2 22
0 9 18
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 3 0
1 U
3835 0 0
2
44799.7 8
0
5 4049~
219 564 396 0 2 22
0 11 19
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 3 0
1 U
3670 0 0
2
44799.7 9
0
5 4049~
219 564 264 0 2 22
0 9 20
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 3 0
1 U
5616 0 0
2
44799.7 10
0
5 4049~
219 564 228 0 2 22
0 11 21
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 3 0
1 U
9323 0 0
2
44799.7 11
0
5 4073~
219 768 576 0 4 22
0 17 13 14 6
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 2 0
1 U
317 0 0
2
44799.7 12
0
5 4073~
219 768 384 0 4 22
0 17 19 18 7
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 1 0
1 U
3108 0 0
2
44799.7 13
0
5 4073~
219 756 204 0 4 22
0 13 21 20 8
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 1 0
1 U
4299 0 0
2
44799.7 14
0
33
5 4 2 0 0 12416 0 13 8 0 0 4
789 756
977 756
977 617
1180 617
3 1 3 0 0 12416 0 7 6 0 0 4
1383 720
1398 720
1398 72
540 72
5 2 4 0 0 4224 0 14 7 0 0 4
789 969
1284 969
1284 729
1337 729
5 1 5 0 0 8320 0 8 7 0 0 4
1230 603
1281 603
1281 711
1337 711
4 3 6 0 0 12416 0 19 8 0 0 4
789 576
925 576
925 608
1180 608
4 0 2 0 0 0 0 8 0 0 1 4
1180 617
1187 617
1187 617
1180 617
4 2 7 0 0 12416 0 20 8 0 0 4
789 384
937 384
937 599
1180 599
1 4 8 0 0 8320 0 8 21 0 0 4
1180 590
965 590
965 204
777 204
0 4 9 0 0 4224 0 0 14 24 0 3
419 432
419 983
744 983
0 3 10 0 0 4224 0 0 14 14 0 3
605 828
605 974
744 974
0 2 11 0 0 8192 0 0 14 16 0 5
246 795
246 941
667 941
667 965
744 965
2 1 12 0 0 4224 0 9 14 0 0 4
588 918
687 918
687 956
744 956
0 1 13 0 0 8192 0 0 9 18 0 3
162 783
162 918
552 918
2 4 10 0 0 0 0 10 13 0 0 4
588 828
709 828
709 770
744 770
0 1 14 0 0 4096 0 0 10 21 0 3
335 585
335 828
552 828
0 3 11 0 0 12416 0 0 13 27 0 6
247 395
246 395
246 796
686 796
686 761
744 761
2 2 15 0 0 4224 0 11 13 0 0 4
588 783
666 783
666 752
744 752
0 1 13 0 0 0 0 0 11 22 0 4
163 576
162 576
162 783
552 783
2 1 16 0 0 8320 0 12 13 0 0 3
585 744
585 743
744 743
0 1 17 0 0 8192 0 0 12 23 0 4
76 567
76 743
549 743
549 744
1 3 14 0 0 4224 0 2 19 0 0 3
335 79
335 585
744 585
0 2 13 0 0 8320 0 0 19 33 0 3
163 195
163 576
744 576
0 1 17 0 0 8320 0 0 19 28 0 3
76 355
76 567
744 567
1 0 9 0 0 0 0 15 0 0 30 3
549 432
419 432
419 260
2 3 18 0 0 4224 0 15 20 0 0 4
585 432
710 432
710 393
744 393
2 2 19 0 0 4224 0 16 20 0 0 4
585 396
686 396
686 384
744 384
0 1 11 0 0 0 0 0 16 32 0 5
246 228
247 228
247 395
549 395
549 396
1 1 17 0 0 0 0 5 20 0 0 4
76 82
76 355
744 355
744 375
2 3 20 0 0 4224 0 17 21 0 0 4
585 264
701 264
701 213
732 213
1 1 9 0 0 0 0 1 17 0 0 3
419 81
419 264
549 264
2 2 21 0 0 4224 0 18 21 0 0 4
585 228
678 228
678 204
732 204
1 1 11 0 0 0 0 3 18 0 0 4
247 82
246 82
246 228
549 228
1 1 13 0 0 0 0 4 21 0 0 3
163 82
163 195
732 195
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
